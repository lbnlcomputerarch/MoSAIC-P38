module full_subtractor_bw8(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a - io_in_b; // @[Arithmetic.scala 42:23]
  wire [9:0] _result_T_2 = _result_T - 9'h0; // @[Arithmetic.scala 42:34]
  wire [8:0] result = _result_T_2[8:0]; // @[Arithmetic.scala 41:22 42:12]
  assign io_out_s = result[7:0]; // @[Arithmetic.scala 43:23]
  assign io_out_c = result[8]; // @[Arithmetic.scala 44:23]
endmodule
module full_adder_bw24(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [23:0] io_out_s,
  output        io_out_c
);
  wire [24:0] _result_T = io_in_a + io_in_b; // @[Arithmetic.scala 27:23]
  wire [25:0] _result_T_1 = {{1'd0}, _result_T}; // @[Arithmetic.scala 27:34]
  wire [24:0] result = _result_T_1[24:0]; // @[Arithmetic.scala 26:22 27:12]
  assign io_out_s = result[23:0]; // @[Arithmetic.scala 28:23]
  assign io_out_c = result[24]; // @[Arithmetic.scala 29:23]
endmodule
module FP_adder_bw32(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] exp_diff_subtractor_io_in_a; // @[FPArithmetic.scala 103:37]
  wire [7:0] exp_diff_subtractor_io_in_b; // @[FPArithmetic.scala 103:37]
  wire [7:0] exp_diff_subtractor_io_out_s; // @[FPArithmetic.scala 103:37]
  wire  exp_diff_subtractor_io_out_c; // @[FPArithmetic.scala 103:37]
  wire [23:0] frac_adder_io_in_a; // @[FPArithmetic.scala 109:28]
  wire [23:0] frac_adder_io_in_b; // @[FPArithmetic.scala 109:28]
  wire [23:0] frac_adder_io_out_s; // @[FPArithmetic.scala 109:28]
  wire  frac_adder_io_out_c; // @[FPArithmetic.scala 109:28]
  wire [7:0] postProcess_exp_diff_subtractor_io_in_a; // @[FPArithmetic.scala 161:49]
  wire [7:0] postProcess_exp_diff_subtractor_io_in_b; // @[FPArithmetic.scala 161:49]
  wire [7:0] postProcess_exp_diff_subtractor_io_out_s; // @[FPArithmetic.scala 161:49]
  wire  postProcess_exp_diff_subtractor_io_out_c; // @[FPArithmetic.scala 161:49]
  wire  sign_wire_0 = io_in_a[31]; // @[FPArithmetic.scala 28:28]
  wire  sign_wire_1 = io_in_b[31]; // @[FPArithmetic.scala 29:28]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 32:64]
  wire [8:0] _GEN_167 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 32:36]
  wire [7:0] _GEN_0 = io_in_a[30:23] < 8'h1 ? 8'h1 : io_in_a[30:23]; // @[FPArithmetic.scala 34:46 35:19 37:19]
  wire [8:0] _GEN_1 = _GEN_167 > _T_2 ? _T_2 : {{1'd0}, _GEN_0}; // @[FPArithmetic.scala 32:71 33:19]
  wire [8:0] _GEN_168 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 39:36]
  wire [7:0] _GEN_2 = io_in_b[30:23] < 8'h1 ? 8'h1 : io_in_b[30:23]; // @[FPArithmetic.scala 41:45 42:19 44:19]
  wire [8:0] _GEN_3 = _GEN_168 > _T_2 ? _T_2 : {{1'd0}, _GEN_2}; // @[FPArithmetic.scala 39:71 40:19]
  wire [22:0] frac_wire_0 = io_in_a[22:0]; // @[FPArithmetic.scala 48:28]
  wire [22:0] frac_wire_1 = io_in_b[22:0]; // @[FPArithmetic.scala 49:28]
  wire [23:0] whole_frac_wire_0 = {1'h1,frac_wire_0}; // @[FPArithmetic.scala 52:31]
  wire [23:0] whole_frac_wire_1 = {1'h1,frac_wire_1}; // @[FPArithmetic.scala 53:31]
  reg  sign_reg_0_0; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_0_1; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_1_0; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_1_1; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_2_0; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_2_1; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_3_0; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_3_1; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_4_0; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_4_1; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_5_0; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_5_1; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_6_0; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_6_1; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_7_0; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_7_1; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_8_0; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_8_1; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_9_0; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_9_1; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_10_0; // @[FPArithmetic.scala 55:27]
  reg  sign_reg_10_1; // @[FPArithmetic.scala 55:27]
  reg [7:0] exp_reg_0_0; // @[FPArithmetic.scala 56:26]
  reg [7:0] exp_reg_0_1; // @[FPArithmetic.scala 56:26]
  reg [7:0] exp_reg_1_0; // @[FPArithmetic.scala 56:26]
  reg [7:0] exp_reg_1_1; // @[FPArithmetic.scala 56:26]
  reg [7:0] exp_reg_2_0; // @[FPArithmetic.scala 56:26]
  reg [7:0] exp_reg_2_1; // @[FPArithmetic.scala 56:26]
  reg [22:0] frac_reg_0_0; // @[FPArithmetic.scala 57:27]
  reg [22:0] frac_reg_0_1; // @[FPArithmetic.scala 57:27]
  reg [22:0] frac_reg_1_0; // @[FPArithmetic.scala 57:27]
  reg [22:0] frac_reg_1_1; // @[FPArithmetic.scala 57:27]
  reg [22:0] frac_reg_2_0; // @[FPArithmetic.scala 57:27]
  reg [22:0] frac_reg_2_1; // @[FPArithmetic.scala 57:27]
  reg [23:0] whole_frac_reg_0_0; // @[FPArithmetic.scala 58:33]
  reg [23:0] whole_frac_reg_0_1; // @[FPArithmetic.scala 58:33]
  reg [23:0] whole_frac_reg_1_0; // @[FPArithmetic.scala 58:33]
  reg [23:0] whole_frac_reg_1_1; // @[FPArithmetic.scala 58:33]
  reg [23:0] whole_frac_reg_2_0; // @[FPArithmetic.scala 58:33]
  reg [23:0] whole_frac_reg_2_1; // @[FPArithmetic.scala 58:33]
  reg [7:0] exp_diff_out_sum_reg_0; // @[FPArithmetic.scala 60:39]
  reg [7:0] exp_diff_out_sum_reg_1; // @[FPArithmetic.scala 60:39]
  reg  exp_diff_out_carry_reg_0; // @[FPArithmetic.scala 61:41]
  reg  exp_diff_out_carry_reg_1; // @[FPArithmetic.scala 61:41]
  reg [23:0] frac_adder_inp_reg_0_0; // @[FPArithmetic.scala 63:37]
  reg [23:0] frac_adder_inp_reg_0_1; // @[FPArithmetic.scala 63:37]
  reg [23:0] frac_adder_inp_reg_1_0; // @[FPArithmetic.scala 63:37]
  reg [23:0] frac_adder_inp_reg_1_1; // @[FPArithmetic.scala 63:37]
  reg  ref_sign_reg_0; // @[FPArithmetic.scala 70:31]
  reg  ref_sign_reg_1; // @[FPArithmetic.scala 70:31]
  reg  ref_sign_reg_2; // @[FPArithmetic.scala 70:31]
  reg  ref_sign_reg_3; // @[FPArithmetic.scala 70:31]
  reg  ref_sign_reg_4; // @[FPArithmetic.scala 70:31]
  reg  ref_sign_reg_5; // @[FPArithmetic.scala 70:31]
  reg  ref_sign_reg_6; // @[FPArithmetic.scala 70:31]
  reg  ref_sign_reg_7; // @[FPArithmetic.scala 70:31]
  reg [22:0] ref_frac_reg_0; // @[FPArithmetic.scala 71:31]
  reg [22:0] ref_frac_reg_1; // @[FPArithmetic.scala 71:31]
  reg [22:0] ref_frac_reg_2; // @[FPArithmetic.scala 71:31]
  reg [22:0] ref_frac_reg_3; // @[FPArithmetic.scala 71:31]
  reg [22:0] ref_frac_reg_4; // @[FPArithmetic.scala 71:31]
  reg [22:0] ref_frac_reg_5; // @[FPArithmetic.scala 71:31]
  reg [22:0] ref_frac_reg_6; // @[FPArithmetic.scala 71:31]
  reg [22:0] ref_frac_reg_7; // @[FPArithmetic.scala 71:31]
  reg [7:0] ref_exp_reg_0; // @[FPArithmetic.scala 72:30]
  reg [7:0] ref_exp_reg_1; // @[FPArithmetic.scala 72:30]
  reg [7:0] ref_exp_reg_2; // @[FPArithmetic.scala 72:30]
  reg [7:0] ref_exp_reg_3; // @[FPArithmetic.scala 72:30]
  reg [7:0] ref_exp_reg_4; // @[FPArithmetic.scala 72:30]
  reg [7:0] ref_exp_reg_5; // @[FPArithmetic.scala 72:30]
  reg [7:0] ref_exp_reg_6; // @[FPArithmetic.scala 72:30]
  reg [7:0] ref_exp_reg_7; // @[FPArithmetic.scala 72:30]
  reg [7:0] ref_exp_diff_reg_0; // @[FPArithmetic.scala 73:35]
  reg [7:0] ref_exp_diff_reg_1; // @[FPArithmetic.scala 73:35]
  reg [7:0] ref_exp_diff_reg_2; // @[FPArithmetic.scala 73:35]
  reg [7:0] ref_exp_diff_reg_3; // @[FPArithmetic.scala 73:35]
  reg [7:0] ref_exp_diff_reg_4; // @[FPArithmetic.scala 73:35]
  reg [7:0] ref_exp_diff_reg_5; // @[FPArithmetic.scala 73:35]
  reg [7:0] ref_exp_diff_reg_6; // @[FPArithmetic.scala 73:35]
  reg [7:0] ref_exp_diff_reg_7; // @[FPArithmetic.scala 73:35]
  reg [23:0] frac_adder_out_sum_reg_0; // @[FPArithmetic.scala 75:41]
  reg [23:0] frac_adder_out_sum_reg_1; // @[FPArithmetic.scala 75:41]
  reg [23:0] frac_adder_out_sum_reg_2; // @[FPArithmetic.scala 75:41]
  reg  frac_adder_out_carry_reg_0; // @[FPArithmetic.scala 76:43]
  reg  new_sign_reg_0; // @[FPArithmetic.scala 82:31]
  reg  new_sign_reg_1; // @[FPArithmetic.scala 82:31]
  reg  new_sign_reg_2; // @[FPArithmetic.scala 82:31]
  reg  new_sign_reg_3; // @[FPArithmetic.scala 82:31]
  reg  new_sign_reg_4; // @[FPArithmetic.scala 82:31]
  reg  new_sign_reg_5; // @[FPArithmetic.scala 82:31]
  reg [22:0] new_frac_reg_0; // @[FPArithmetic.scala 83:31]
  reg [7:0] new_exp_reg_0; // @[FPArithmetic.scala 84:30]
  reg  noPostProcess_reg_0; // @[FPArithmetic.scala 89:36]
  reg  noPostProcess_reg_1; // @[FPArithmetic.scala 89:36]
  reg  noPostProcess_reg_2; // @[FPArithmetic.scala 89:36]
  reg  noPostProcess_reg_3; // @[FPArithmetic.scala 89:36]
  reg  noPostProcess_reg_4; // @[FPArithmetic.scala 89:36]
  reg  postProcessInstruction_reg_0; // @[FPArithmetic.scala 90:45]
  reg  postProcessInstruction_reg_1; // @[FPArithmetic.scala 90:45]
  reg  postProcessInstruction_reg_2; // @[FPArithmetic.scala 90:45]
  reg  postProcessInstruction_reg_3; // @[FPArithmetic.scala 90:45]
  reg  postProcessInstruction_reg_4; // @[FPArithmetic.scala 90:45]
  reg [23:0] ref_frac_adder_sum_reg_0; // @[FPArithmetic.scala 92:41]
  reg [23:0] ref_frac_adder_sum_reg_1; // @[FPArithmetic.scala 92:41]
  reg [23:0] ref_frac_adder_sum_reg_2; // @[FPArithmetic.scala 92:41]
  reg [5:0] leadingOne_reg_0; // @[FPArithmetic.scala 94:33]
  reg [5:0] leadingOne_reg_1; // @[FPArithmetic.scala 94:33]
  reg [31:0] input_a_reg_0; // @[FPArithmetic.scala 96:30]
  reg [31:0] input_a_reg_1; // @[FPArithmetic.scala 96:30]
  reg [31:0] input_a_reg_2; // @[FPArithmetic.scala 96:30]
  reg [31:0] input_a_reg_3; // @[FPArithmetic.scala 96:30]
  reg [31:0] input_a_reg_4; // @[FPArithmetic.scala 96:30]
  reg [31:0] input_a_reg_5; // @[FPArithmetic.scala 96:30]
  reg [31:0] input_a_reg_6; // @[FPArithmetic.scala 96:30]
  reg [31:0] input_a_reg_7; // @[FPArithmetic.scala 96:30]
  reg [31:0] input_a_reg_8; // @[FPArithmetic.scala 96:30]
  reg [31:0] input_a_reg_9; // @[FPArithmetic.scala 96:30]
  reg [31:0] input_a_reg_10; // @[FPArithmetic.scala 96:30]
  reg [31:0] input_b_reg_0; // @[FPArithmetic.scala 97:30]
  reg [31:0] input_b_reg_1; // @[FPArithmetic.scala 97:30]
  reg [31:0] input_b_reg_2; // @[FPArithmetic.scala 97:30]
  reg [31:0] input_b_reg_3; // @[FPArithmetic.scala 97:30]
  reg [31:0] input_b_reg_4; // @[FPArithmetic.scala 97:30]
  reg [31:0] input_b_reg_5; // @[FPArithmetic.scala 97:30]
  reg [31:0] input_b_reg_6; // @[FPArithmetic.scala 97:30]
  reg [31:0] input_b_reg_7; // @[FPArithmetic.scala 97:30]
  reg [31:0] input_b_reg_8; // @[FPArithmetic.scala 97:30]
  reg [31:0] input_b_reg_9; // @[FPArithmetic.scala 97:30]
  reg [31:0] input_b_reg_10; // @[FPArithmetic.scala 97:30]
  reg [7:0] postProcess_exp_diff_out_sum_reg_0; // @[FPArithmetic.scala 99:51]
  reg  postProcess_exp_diff_out_carry_reg_0; // @[FPArithmetic.scala 100:53]
  reg [7:0] cmpl_subber_out_s_reg_0; // @[FPArithmetic.scala 114:40]
  wire [7:0] _cmpl_subber_out_s_reg_0_T = ~exp_diff_out_sum_reg_0; // @[FPArithmetic.scala 116:41]
  wire [7:0] _cmpl_subber_out_s_reg_0_T_2 = 8'h1 + _cmpl_subber_out_s_reg_0_T; // @[FPArithmetic.scala 116:39]
  wire [23:0] _frac_adder_inp_wire_0_T = whole_frac_reg_2_0 >> cmpl_subber_out_s_reg_0; // @[FPArithmetic.scala 124:54]
  wire [23:0] _frac_adder_inp_wire_1_T = whole_frac_reg_2_1 >> exp_diff_out_sum_reg_1; // @[FPArithmetic.scala 132:54]
  reg [23:0] cmpl_frac_adder_inp_reg_0_0; // @[FPArithmetic.scala 135:42]
  reg [23:0] cmpl_frac_adder_inp_reg_0_1; // @[FPArithmetic.scala 135:42]
  wire [23:0] _cmpl_frac_adder_inp_reg_0_0_T = ~frac_adder_inp_reg_0_0; // @[FPArithmetic.scala 137:46]
  wire [23:0] _cmpl_frac_adder_inp_reg_0_0_T_2 = 24'h1 + _cmpl_frac_adder_inp_reg_0_0_T; // @[FPArithmetic.scala 137:44]
  wire [23:0] _cmpl_frac_adder_inp_reg_0_1_T = ~frac_adder_inp_reg_0_1; // @[FPArithmetic.scala 138:46]
  wire [23:0] _cmpl_frac_adder_inp_reg_0_1_T_2 = 24'h1 + _cmpl_frac_adder_inp_reg_0_1_T; // @[FPArithmetic.scala 138:44]
  wire [1:0] _frac_adder_io_in_a_T = {sign_reg_4_1,sign_reg_4_0}; // @[FPArithmetic.scala 141:43]
  wire  _new_sign_wire_T = ~frac_adder_out_carry_reg_0; // @[FPArithmetic.scala 144:23]
  wire  new_sign_wire = ~frac_adder_out_carry_reg_0 & (sign_reg_5_0 | sign_reg_5_1) | sign_reg_5_0 & sign_reg_5_1; // @[FPArithmetic.scala 144:89]
  wire  _noPostProcess_wire_T_5 = sign_reg_5_0 ^ sign_reg_5_1; // @[FPArithmetic.scala 148:148]
  wire  noPostProcess_wire = _new_sign_wire_T & ~frac_adder_out_sum_reg_0[23] | _new_sign_wire_T & ~(sign_reg_5_0 ^
    sign_reg_5_1) | frac_adder_out_carry_reg_0 & frac_adder_out_sum_reg_0[23] & (sign_reg_5_0 ^ sign_reg_5_1); // @[FPArithmetic.scala 148:167]
  wire  postProcessInstruction_wire = _new_sign_wire_T | _noPostProcess_wire_T_5; // @[FPArithmetic.scala 149:67]
  reg [23:0] cmpl_frac_adder_out_sum_reg_0; // @[FPArithmetic.scala 151:46]
  wire [23:0] _cmpl_frac_adder_out_sum_reg_0_T = ~frac_adder_out_sum_reg_1; // @[FPArithmetic.scala 153:47]
  wire [23:0] _cmpl_frac_adder_out_sum_reg_0_T_2 = 24'h1 + _cmpl_frac_adder_out_sum_reg_0_T; // @[FPArithmetic.scala 153:45]
  wire [1:0] _ref_frac_adder_sum_wire_T = {sign_reg_7_1,sign_reg_7_0}; // @[FPArithmetic.scala 157:67]
  wire [1:0] _leadingOne_wire_T_25 = ref_frac_adder_sum_reg_0[2] ? 2'h2 : {{1'd0}, ref_frac_adder_sum_reg_0[1]}; // @[FPArithmetic.scala 160:81]
  wire [1:0] _leadingOne_wire_T_26 = ref_frac_adder_sum_reg_0[3] ? 2'h3 : _leadingOne_wire_T_25; // @[FPArithmetic.scala 160:81]
  wire [2:0] _leadingOne_wire_T_27 = ref_frac_adder_sum_reg_0[4] ? 3'h4 : {{1'd0}, _leadingOne_wire_T_26}; // @[FPArithmetic.scala 160:81]
  wire [2:0] _leadingOne_wire_T_28 = ref_frac_adder_sum_reg_0[5] ? 3'h5 : _leadingOne_wire_T_27; // @[FPArithmetic.scala 160:81]
  wire [2:0] _leadingOne_wire_T_29 = ref_frac_adder_sum_reg_0[6] ? 3'h6 : _leadingOne_wire_T_28; // @[FPArithmetic.scala 160:81]
  wire [2:0] _leadingOne_wire_T_30 = ref_frac_adder_sum_reg_0[7] ? 3'h7 : _leadingOne_wire_T_29; // @[FPArithmetic.scala 160:81]
  wire [3:0] _leadingOne_wire_T_31 = ref_frac_adder_sum_reg_0[8] ? 4'h8 : {{1'd0}, _leadingOne_wire_T_30}; // @[FPArithmetic.scala 160:81]
  wire [3:0] _leadingOne_wire_T_32 = ref_frac_adder_sum_reg_0[9] ? 4'h9 : _leadingOne_wire_T_31; // @[FPArithmetic.scala 160:81]
  wire [3:0] _leadingOne_wire_T_33 = ref_frac_adder_sum_reg_0[10] ? 4'ha : _leadingOne_wire_T_32; // @[FPArithmetic.scala 160:81]
  wire [3:0] _leadingOne_wire_T_34 = ref_frac_adder_sum_reg_0[11] ? 4'hb : _leadingOne_wire_T_33; // @[FPArithmetic.scala 160:81]
  wire [3:0] _leadingOne_wire_T_35 = ref_frac_adder_sum_reg_0[12] ? 4'hc : _leadingOne_wire_T_34; // @[FPArithmetic.scala 160:81]
  wire [3:0] _leadingOne_wire_T_36 = ref_frac_adder_sum_reg_0[13] ? 4'hd : _leadingOne_wire_T_35; // @[FPArithmetic.scala 160:81]
  wire [3:0] _leadingOne_wire_T_37 = ref_frac_adder_sum_reg_0[14] ? 4'he : _leadingOne_wire_T_36; // @[FPArithmetic.scala 160:81]
  wire [3:0] _leadingOne_wire_T_38 = ref_frac_adder_sum_reg_0[15] ? 4'hf : _leadingOne_wire_T_37; // @[FPArithmetic.scala 160:81]
  wire [4:0] _leadingOne_wire_T_39 = ref_frac_adder_sum_reg_0[16] ? 5'h10 : {{1'd0}, _leadingOne_wire_T_38}; // @[FPArithmetic.scala 160:81]
  wire [4:0] _leadingOne_wire_T_40 = ref_frac_adder_sum_reg_0[17] ? 5'h11 : _leadingOne_wire_T_39; // @[FPArithmetic.scala 160:81]
  wire [4:0] _leadingOne_wire_T_41 = ref_frac_adder_sum_reg_0[18] ? 5'h12 : _leadingOne_wire_T_40; // @[FPArithmetic.scala 160:81]
  wire [4:0] _leadingOne_wire_T_42 = ref_frac_adder_sum_reg_0[19] ? 5'h13 : _leadingOne_wire_T_41; // @[FPArithmetic.scala 160:81]
  wire [4:0] _leadingOne_wire_T_43 = ref_frac_adder_sum_reg_0[20] ? 5'h14 : _leadingOne_wire_T_42; // @[FPArithmetic.scala 160:81]
  wire [4:0] _leadingOne_wire_T_44 = ref_frac_adder_sum_reg_0[21] ? 5'h15 : _leadingOne_wire_T_43; // @[FPArithmetic.scala 160:81]
  wire [4:0] _leadingOne_wire_T_45 = ref_frac_adder_sum_reg_0[22] ? 5'h16 : _leadingOne_wire_T_44; // @[FPArithmetic.scala 160:81]
  wire [4:0] _leadingOne_wire_T_46 = ref_frac_adder_sum_reg_0[23] ? 5'h17 : _leadingOne_wire_T_45; // @[FPArithmetic.scala 160:81]
  wire [5:0] leadingOne_wire = _leadingOne_wire_T_46 + 5'h1; // @[FPArithmetic.scala 160:88]
  wire [5:0] _postProcess_exp_diff_subtractor_io_in_b_T_1 = 6'h18 - leadingOne_reg_0; // @[FPArithmetic.scala 163:66]
  wire [7:0] exp_wire_0 = _GEN_1[7:0]; // @[FPArithmetic.scala 30:24]
  wire [7:0] exp_wire_1 = _GEN_3[7:0]; // @[FPArithmetic.scala 30:24]
  reg [31:0] output_sum_reg; // @[FPArithmetic.scala 221:33]
  wire [8:0] _GEN_169 = {{1'd0}, ref_exp_reg_7}; // @[FPArithmetic.scala 238:29]
  wire [23:0] _new_frac_reg_0_T_2 = 24'h800000 - 24'h1; // @[FPArithmetic.scala 240:56]
  wire [7:0] _new_exp_reg_0_T_3 = ref_exp_reg_7 + 8'h1; // @[FPArithmetic.scala 242:44]
  wire [8:0] _GEN_142 = _GEN_169 == _T_2 ? _T_2 : {{1'd0}, _new_exp_reg_0_T_3}; // @[FPArithmetic.scala 238:66 239:26 242:26]
  wire [23:0] _GEN_143 = _GEN_169 == _T_2 ? _new_frac_reg_0_T_2 : {{1'd0}, ref_frac_adder_sum_reg_2[23:1]}; // @[FPArithmetic.scala 238:66 240:27 243:27]
  wire [5:0] _new_frac_reg_0_T_6 = 6'h18 - leadingOne_reg_1; // @[FPArithmetic.scala 256:96]
  wire [85:0] _GEN_5 = {{63'd0}, ref_frac_adder_sum_reg_2[22:0]}; // @[FPArithmetic.scala 256:75]
  wire [85:0] _new_frac_reg_0_T_7 = _GEN_5 << _new_frac_reg_0_T_6; // @[FPArithmetic.scala 256:75]
  wire [7:0] _GEN_144 = postProcess_exp_diff_out_carry_reg_0 ? 8'h1 : postProcess_exp_diff_out_sum_reg_0; // @[FPArithmetic.scala 251:63 252:28 255:28]
  wire [85:0] _GEN_145 = postProcess_exp_diff_out_carry_reg_0 ? 86'h0 : _new_frac_reg_0_T_7; // @[FPArithmetic.scala 251:63 253:29 256:29]
  wire [7:0] _GEN_146 = leadingOne_reg_1 == 6'h1 & ref_frac_adder_sum_reg_2 == 24'h0 & ((sign_reg_10_0 ^ sign_reg_10_1)
     & input_a_reg_10[30:0] == input_b_reg_10[30:0]) ? 8'h0 : _GEN_144; // @[FPArithmetic.scala 247:190 248:26]
  wire [85:0] _GEN_147 = leadingOne_reg_1 == 6'h1 & ref_frac_adder_sum_reg_2 == 24'h0 & ((sign_reg_10_0 ^ sign_reg_10_1)
     & input_a_reg_10[30:0] == input_b_reg_10[30:0]) ? 86'h0 : _GEN_145; // @[FPArithmetic.scala 247:190 249:27]
  wire  _GEN_148 = postProcessInstruction_reg_4 ? new_sign_reg_4 : new_sign_reg_5; // @[FPArithmetic.scala 245:57 246:25 82:31]
  wire [7:0] _GEN_149 = postProcessInstruction_reg_4 ? _GEN_146 : new_exp_reg_0; // @[FPArithmetic.scala 245:57 84:30]
  wire [85:0] _GEN_150 = postProcessInstruction_reg_4 ? _GEN_147 : {{63'd0}, new_frac_reg_0}; // @[FPArithmetic.scala 245:57 83:31]
  wire  _GEN_151 = ~postProcessInstruction_reg_4 ? new_sign_reg_4 : _GEN_148; // @[FPArithmetic.scala 236:57 237:25]
  wire [8:0] _GEN_152 = ~postProcessInstruction_reg_4 ? _GEN_142 : {{1'd0}, _GEN_149}; // @[FPArithmetic.scala 236:57]
  wire [85:0] _GEN_153 = ~postProcessInstruction_reg_4 ? {{62'd0}, _GEN_143} : _GEN_150; // @[FPArithmetic.scala 236:57]
  wire  _GEN_154 = noPostProcess_reg_4 ? new_sign_reg_4 : _GEN_151; // @[FPArithmetic.scala 232:48 233:25]
  wire [8:0] _GEN_155 = noPostProcess_reg_4 ? {{1'd0}, ref_exp_reg_7} : _GEN_152; // @[FPArithmetic.scala 232:48 234:24]
  wire [85:0] _GEN_156 = noPostProcess_reg_4 ? {{63'd0}, ref_frac_adder_sum_reg_2[22:0]} : _GEN_153; // @[FPArithmetic.scala 232:48 235:25]
  wire [85:0] _GEN_158 = ref_exp_diff_reg_7 >= 8'h17 ? {{63'd0}, ref_frac_reg_7} : _GEN_156; // @[FPArithmetic.scala 228:53 230:25]
  wire [8:0] _GEN_159 = ref_exp_diff_reg_7 >= 8'h17 ? {{1'd0}, ref_exp_reg_7} : _GEN_155; // @[FPArithmetic.scala 228:53 231:24]
  wire [8:0] _GEN_161 = input_a_reg_10[30:0] == 31'h0 & input_b_reg_10[30:0] == 31'h0 ? 9'h0 : _GEN_159; // @[FPArithmetic.scala 224:86 226:24]
  wire [85:0] _GEN_162 = input_a_reg_10[30:0] == 31'h0 & input_b_reg_10[30:0] == 31'h0 ? 86'h0 : _GEN_158; // @[FPArithmetic.scala 224:86 227:25]
  wire [31:0] _output_sum_reg_T_1 = {new_sign_reg_5,new_exp_reg_0,new_frac_reg_0}; // @[FPArithmetic.scala 260:59]
  wire [8:0] _GEN_164 = io_in_en ? _GEN_161 : {{1'd0}, new_exp_reg_0}; // @[FPArithmetic.scala 223:20 84:30]
  wire [85:0] _GEN_165 = io_in_en ? _GEN_162 : {{63'd0}, new_frac_reg_0}; // @[FPArithmetic.scala 223:20 83:31]
  wire [85:0] _GEN_170 = reset ? 86'h0 : _GEN_165; // @[FPArithmetic.scala 83:{31,31}]
  wire [8:0] _GEN_171 = reset ? 9'h0 : _GEN_164; // @[FPArithmetic.scala 84:{30,30}]
  full_subtractor_bw8 exp_diff_subtractor ( // @[FPArithmetic.scala 103:37]
    .io_in_a(exp_diff_subtractor_io_in_a),
    .io_in_b(exp_diff_subtractor_io_in_b),
    .io_out_s(exp_diff_subtractor_io_out_s),
    .io_out_c(exp_diff_subtractor_io_out_c)
  );
  full_adder_bw24 frac_adder ( // @[FPArithmetic.scala 109:28]
    .io_in_a(frac_adder_io_in_a),
    .io_in_b(frac_adder_io_in_b),
    .io_out_s(frac_adder_io_out_s),
    .io_out_c(frac_adder_io_out_c)
  );
  full_subtractor_bw8 postProcess_exp_diff_subtractor ( // @[FPArithmetic.scala 161:49]
    .io_in_a(postProcess_exp_diff_subtractor_io_in_a),
    .io_in_b(postProcess_exp_diff_subtractor_io_in_b),
    .io_out_s(postProcess_exp_diff_subtractor_io_out_s),
    .io_out_c(postProcess_exp_diff_subtractor_io_out_c)
  );
  assign io_out_s = output_sum_reg; // @[FPArithmetic.scala 222:14]
  assign exp_diff_subtractor_io_in_a = exp_reg_0_0; // @[FPArithmetic.scala 104:33]
  assign exp_diff_subtractor_io_in_b = exp_reg_0_1; // @[FPArithmetic.scala 105:33]
  assign frac_adder_io_in_a = _frac_adder_io_in_a_T == 2'h1 ? cmpl_frac_adder_inp_reg_0_0 : frac_adder_inp_reg_1_0; // @[FPArithmetic.scala 141:30]
  assign frac_adder_io_in_b = _frac_adder_io_in_a_T == 2'h2 ? cmpl_frac_adder_inp_reg_0_1 : frac_adder_inp_reg_1_1; // @[FPArithmetic.scala 142:30]
  assign postProcess_exp_diff_subtractor_io_in_a = ref_exp_reg_6; // @[FPArithmetic.scala 162:45]
  assign postProcess_exp_diff_subtractor_io_in_b = {{2'd0}, _postProcess_exp_diff_subtractor_io_in_b_T_1}; // @[FPArithmetic.scala 163:45]
  always @(posedge clock) begin
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_0_0 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_0_0 <= sign_wire_0; // @[FPArithmetic.scala 169:19]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_0_1 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_0_1 <= sign_wire_1; // @[FPArithmetic.scala 169:19]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_1_0 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_1_0 <= sign_reg_0_0; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_1_1 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_1_1 <= sign_reg_0_1; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_2_0 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_2_0 <= sign_reg_1_0; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_2_1 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_2_1 <= sign_reg_1_1; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_3_0 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_3_0 <= sign_reg_2_0; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_3_1 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_3_1 <= sign_reg_2_1; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_4_0 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_4_0 <= sign_reg_3_0; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_4_1 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_4_1 <= sign_reg_3_1; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_5_0 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_5_0 <= sign_reg_4_0; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_5_1 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_5_1 <= sign_reg_4_1; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_6_0 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_6_0 <= sign_reg_5_0; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_6_1 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_6_1 <= sign_reg_5_1; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_7_0 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_7_0 <= sign_reg_6_0; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_7_1 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_7_1 <= sign_reg_6_1; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_8_0 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_8_0 <= sign_reg_7_0; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_8_1 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_8_1 <= sign_reg_7_1; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_9_0 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_9_0 <= sign_reg_8_0; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_9_1 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_9_1 <= sign_reg_8_1; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_10_0 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_10_0 <= sign_reg_9_0; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 55:27]
      sign_reg_10_1 <= 1'h0; // @[FPArithmetic.scala 55:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      sign_reg_10_1 <= sign_reg_9_1; // @[FPArithmetic.scala 191:23]
    end
    if (reset) begin // @[FPArithmetic.scala 56:26]
      exp_reg_0_0 <= 8'h0; // @[FPArithmetic.scala 56:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      exp_reg_0_0 <= exp_wire_0; // @[FPArithmetic.scala 170:18]
    end
    if (reset) begin // @[FPArithmetic.scala 56:26]
      exp_reg_0_1 <= 8'h0; // @[FPArithmetic.scala 56:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      exp_reg_0_1 <= exp_wire_1; // @[FPArithmetic.scala 170:18]
    end
    if (reset) begin // @[FPArithmetic.scala 56:26]
      exp_reg_1_0 <= 8'h0; // @[FPArithmetic.scala 56:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      exp_reg_1_0 <= exp_reg_0_0; // @[FPArithmetic.scala 209:22]
    end
    if (reset) begin // @[FPArithmetic.scala 56:26]
      exp_reg_1_1 <= 8'h0; // @[FPArithmetic.scala 56:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      exp_reg_1_1 <= exp_reg_0_1; // @[FPArithmetic.scala 209:22]
    end
    if (reset) begin // @[FPArithmetic.scala 56:26]
      exp_reg_2_0 <= 8'h0; // @[FPArithmetic.scala 56:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      exp_reg_2_0 <= exp_reg_1_0; // @[FPArithmetic.scala 209:22]
    end
    if (reset) begin // @[FPArithmetic.scala 56:26]
      exp_reg_2_1 <= 8'h0; // @[FPArithmetic.scala 56:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      exp_reg_2_1 <= exp_reg_1_1; // @[FPArithmetic.scala 209:22]
    end
    if (reset) begin // @[FPArithmetic.scala 57:27]
      frac_reg_0_0 <= 23'h0; // @[FPArithmetic.scala 57:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      frac_reg_0_0 <= frac_wire_0; // @[FPArithmetic.scala 171:19]
    end
    if (reset) begin // @[FPArithmetic.scala 57:27]
      frac_reg_0_1 <= 23'h0; // @[FPArithmetic.scala 57:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      frac_reg_0_1 <= frac_wire_1; // @[FPArithmetic.scala 171:19]
    end
    if (reset) begin // @[FPArithmetic.scala 57:27]
      frac_reg_1_0 <= 23'h0; // @[FPArithmetic.scala 57:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      frac_reg_1_0 <= frac_reg_0_0; // @[FPArithmetic.scala 210:23]
    end
    if (reset) begin // @[FPArithmetic.scala 57:27]
      frac_reg_1_1 <= 23'h0; // @[FPArithmetic.scala 57:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      frac_reg_1_1 <= frac_reg_0_1; // @[FPArithmetic.scala 210:23]
    end
    if (reset) begin // @[FPArithmetic.scala 57:27]
      frac_reg_2_0 <= 23'h0; // @[FPArithmetic.scala 57:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      frac_reg_2_0 <= frac_reg_1_0; // @[FPArithmetic.scala 210:23]
    end
    if (reset) begin // @[FPArithmetic.scala 57:27]
      frac_reg_2_1 <= 23'h0; // @[FPArithmetic.scala 57:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      frac_reg_2_1 <= frac_reg_1_1; // @[FPArithmetic.scala 210:23]
    end
    if (reset) begin // @[FPArithmetic.scala 58:33]
      whole_frac_reg_0_0 <= 24'h0; // @[FPArithmetic.scala 58:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      whole_frac_reg_0_0 <= whole_frac_wire_0; // @[FPArithmetic.scala 172:25]
    end
    if (reset) begin // @[FPArithmetic.scala 58:33]
      whole_frac_reg_0_1 <= 24'h0; // @[FPArithmetic.scala 58:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      whole_frac_reg_0_1 <= whole_frac_wire_1; // @[FPArithmetic.scala 172:25]
    end
    if (reset) begin // @[FPArithmetic.scala 58:33]
      whole_frac_reg_1_0 <= 24'h0; // @[FPArithmetic.scala 58:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      whole_frac_reg_1_0 <= whole_frac_reg_0_0; // @[FPArithmetic.scala 211:29]
    end
    if (reset) begin // @[FPArithmetic.scala 58:33]
      whole_frac_reg_1_1 <= 24'h0; // @[FPArithmetic.scala 58:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      whole_frac_reg_1_1 <= whole_frac_reg_0_1; // @[FPArithmetic.scala 211:29]
    end
    if (reset) begin // @[FPArithmetic.scala 58:33]
      whole_frac_reg_2_0 <= 24'h0; // @[FPArithmetic.scala 58:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      whole_frac_reg_2_0 <= whole_frac_reg_1_0; // @[FPArithmetic.scala 211:29]
    end
    if (reset) begin // @[FPArithmetic.scala 58:33]
      whole_frac_reg_2_1 <= 24'h0; // @[FPArithmetic.scala 58:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      whole_frac_reg_2_1 <= whole_frac_reg_1_1; // @[FPArithmetic.scala 211:29]
    end
    if (reset) begin // @[FPArithmetic.scala 60:39]
      exp_diff_out_sum_reg_0 <= 8'h0; // @[FPArithmetic.scala 60:39]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      exp_diff_out_sum_reg_0 <= exp_diff_subtractor_io_out_s; // @[FPArithmetic.scala 173:31]
    end
    if (reset) begin // @[FPArithmetic.scala 60:39]
      exp_diff_out_sum_reg_1 <= 8'h0; // @[FPArithmetic.scala 60:39]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      exp_diff_out_sum_reg_1 <= exp_diff_out_sum_reg_0; // @[FPArithmetic.scala 214:35]
    end
    if (reset) begin // @[FPArithmetic.scala 61:41]
      exp_diff_out_carry_reg_0 <= 1'h0; // @[FPArithmetic.scala 61:41]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      exp_diff_out_carry_reg_0 <= exp_diff_subtractor_io_out_c; // @[FPArithmetic.scala 174:33]
    end
    if (reset) begin // @[FPArithmetic.scala 61:41]
      exp_diff_out_carry_reg_1 <= 1'h0; // @[FPArithmetic.scala 61:41]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      exp_diff_out_carry_reg_1 <= exp_diff_out_carry_reg_0; // @[FPArithmetic.scala 215:37]
    end
    if (reset) begin // @[FPArithmetic.scala 63:37]
      frac_adder_inp_reg_0_0 <= 24'h0; // @[FPArithmetic.scala 63:37]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      if (exp_diff_out_carry_reg_1) begin // @[FPArithmetic.scala 119:45]
        frac_adder_inp_reg_0_0 <= _frac_adder_inp_wire_0_T; // @[FPArithmetic.scala 124:30]
      end else begin
        frac_adder_inp_reg_0_0 <= whole_frac_reg_2_0; // @[FPArithmetic.scala 131:30]
      end
    end
    if (reset) begin // @[FPArithmetic.scala 63:37]
      frac_adder_inp_reg_0_1 <= 24'h0; // @[FPArithmetic.scala 63:37]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      if (exp_diff_out_carry_reg_1) begin // @[FPArithmetic.scala 119:45]
        frac_adder_inp_reg_0_1 <= whole_frac_reg_2_1; // @[FPArithmetic.scala 125:30]
      end else begin
        frac_adder_inp_reg_0_1 <= _frac_adder_inp_wire_1_T; // @[FPArithmetic.scala 132:30]
      end
    end
    if (reset) begin // @[FPArithmetic.scala 63:37]
      frac_adder_inp_reg_1_0 <= 24'h0; // @[FPArithmetic.scala 63:37]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      frac_adder_inp_reg_1_0 <= frac_adder_inp_reg_0_0; // @[FPArithmetic.scala 217:33]
    end
    if (reset) begin // @[FPArithmetic.scala 63:37]
      frac_adder_inp_reg_1_1 <= 24'h0; // @[FPArithmetic.scala 63:37]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      frac_adder_inp_reg_1_1 <= frac_adder_inp_reg_0_1; // @[FPArithmetic.scala 217:33]
    end
    if (reset) begin // @[FPArithmetic.scala 70:31]
      ref_sign_reg_0 <= 1'h0; // @[FPArithmetic.scala 70:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      if (exp_diff_out_carry_reg_1) begin // @[FPArithmetic.scala 119:45]
        ref_sign_reg_0 <= sign_reg_2_1; // @[FPArithmetic.scala 122:21]
      end else begin
        ref_sign_reg_0 <= sign_reg_2_0; // @[FPArithmetic.scala 129:21]
      end
    end
    if (reset) begin // @[FPArithmetic.scala 70:31]
      ref_sign_reg_1 <= 1'h0; // @[FPArithmetic.scala 70:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_sign_reg_1 <= ref_sign_reg_0; // @[FPArithmetic.scala 196:27]
    end
    if (reset) begin // @[FPArithmetic.scala 70:31]
      ref_sign_reg_2 <= 1'h0; // @[FPArithmetic.scala 70:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_sign_reg_2 <= ref_sign_reg_1; // @[FPArithmetic.scala 196:27]
    end
    if (reset) begin // @[FPArithmetic.scala 70:31]
      ref_sign_reg_3 <= 1'h0; // @[FPArithmetic.scala 70:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_sign_reg_3 <= ref_sign_reg_2; // @[FPArithmetic.scala 196:27]
    end
    if (reset) begin // @[FPArithmetic.scala 70:31]
      ref_sign_reg_4 <= 1'h0; // @[FPArithmetic.scala 70:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_sign_reg_4 <= ref_sign_reg_3; // @[FPArithmetic.scala 196:27]
    end
    if (reset) begin // @[FPArithmetic.scala 70:31]
      ref_sign_reg_5 <= 1'h0; // @[FPArithmetic.scala 70:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_sign_reg_5 <= ref_sign_reg_4; // @[FPArithmetic.scala 196:27]
    end
    if (reset) begin // @[FPArithmetic.scala 70:31]
      ref_sign_reg_6 <= 1'h0; // @[FPArithmetic.scala 70:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_sign_reg_6 <= ref_sign_reg_5; // @[FPArithmetic.scala 196:27]
    end
    if (reset) begin // @[FPArithmetic.scala 70:31]
      ref_sign_reg_7 <= 1'h0; // @[FPArithmetic.scala 70:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_sign_reg_7 <= ref_sign_reg_6; // @[FPArithmetic.scala 196:27]
    end
    if (reset) begin // @[FPArithmetic.scala 71:31]
      ref_frac_reg_0 <= 23'h0; // @[FPArithmetic.scala 71:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      if (exp_diff_out_carry_reg_1) begin // @[FPArithmetic.scala 119:45]
        ref_frac_reg_0 <= frac_reg_2_1; // @[FPArithmetic.scala 123:21]
      end else begin
        ref_frac_reg_0 <= frac_reg_2_0; // @[FPArithmetic.scala 130:21]
      end
    end
    if (reset) begin // @[FPArithmetic.scala 71:31]
      ref_frac_reg_1 <= 23'h0; // @[FPArithmetic.scala 71:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_frac_reg_1 <= ref_frac_reg_0; // @[FPArithmetic.scala 197:27]
    end
    if (reset) begin // @[FPArithmetic.scala 71:31]
      ref_frac_reg_2 <= 23'h0; // @[FPArithmetic.scala 71:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_frac_reg_2 <= ref_frac_reg_1; // @[FPArithmetic.scala 197:27]
    end
    if (reset) begin // @[FPArithmetic.scala 71:31]
      ref_frac_reg_3 <= 23'h0; // @[FPArithmetic.scala 71:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_frac_reg_3 <= ref_frac_reg_2; // @[FPArithmetic.scala 197:27]
    end
    if (reset) begin // @[FPArithmetic.scala 71:31]
      ref_frac_reg_4 <= 23'h0; // @[FPArithmetic.scala 71:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_frac_reg_4 <= ref_frac_reg_3; // @[FPArithmetic.scala 197:27]
    end
    if (reset) begin // @[FPArithmetic.scala 71:31]
      ref_frac_reg_5 <= 23'h0; // @[FPArithmetic.scala 71:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_frac_reg_5 <= ref_frac_reg_4; // @[FPArithmetic.scala 197:27]
    end
    if (reset) begin // @[FPArithmetic.scala 71:31]
      ref_frac_reg_6 <= 23'h0; // @[FPArithmetic.scala 71:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_frac_reg_6 <= ref_frac_reg_5; // @[FPArithmetic.scala 197:27]
    end
    if (reset) begin // @[FPArithmetic.scala 71:31]
      ref_frac_reg_7 <= 23'h0; // @[FPArithmetic.scala 71:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_frac_reg_7 <= ref_frac_reg_6; // @[FPArithmetic.scala 197:27]
    end
    if (reset) begin // @[FPArithmetic.scala 72:30]
      ref_exp_reg_0 <= 8'h0; // @[FPArithmetic.scala 72:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      if (exp_diff_out_carry_reg_1) begin // @[FPArithmetic.scala 119:45]
        ref_exp_reg_0 <= exp_reg_2_1; // @[FPArithmetic.scala 120:20]
      end else begin
        ref_exp_reg_0 <= exp_reg_2_0; // @[FPArithmetic.scala 127:20]
      end
    end
    if (reset) begin // @[FPArithmetic.scala 72:30]
      ref_exp_reg_1 <= 8'h0; // @[FPArithmetic.scala 72:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_reg_1 <= ref_exp_reg_0; // @[FPArithmetic.scala 198:26]
    end
    if (reset) begin // @[FPArithmetic.scala 72:30]
      ref_exp_reg_2 <= 8'h0; // @[FPArithmetic.scala 72:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_reg_2 <= ref_exp_reg_1; // @[FPArithmetic.scala 198:26]
    end
    if (reset) begin // @[FPArithmetic.scala 72:30]
      ref_exp_reg_3 <= 8'h0; // @[FPArithmetic.scala 72:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_reg_3 <= ref_exp_reg_2; // @[FPArithmetic.scala 198:26]
    end
    if (reset) begin // @[FPArithmetic.scala 72:30]
      ref_exp_reg_4 <= 8'h0; // @[FPArithmetic.scala 72:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_reg_4 <= ref_exp_reg_3; // @[FPArithmetic.scala 198:26]
    end
    if (reset) begin // @[FPArithmetic.scala 72:30]
      ref_exp_reg_5 <= 8'h0; // @[FPArithmetic.scala 72:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_reg_5 <= ref_exp_reg_4; // @[FPArithmetic.scala 198:26]
    end
    if (reset) begin // @[FPArithmetic.scala 72:30]
      ref_exp_reg_6 <= 8'h0; // @[FPArithmetic.scala 72:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_reg_6 <= ref_exp_reg_5; // @[FPArithmetic.scala 198:26]
    end
    if (reset) begin // @[FPArithmetic.scala 72:30]
      ref_exp_reg_7 <= 8'h0; // @[FPArithmetic.scala 72:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_reg_7 <= ref_exp_reg_6; // @[FPArithmetic.scala 198:26]
    end
    if (reset) begin // @[FPArithmetic.scala 73:35]
      ref_exp_diff_reg_0 <= 8'h0; // @[FPArithmetic.scala 73:35]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      if (exp_diff_out_carry_reg_1) begin // @[FPArithmetic.scala 119:45]
        ref_exp_diff_reg_0 <= cmpl_subber_out_s_reg_0; // @[FPArithmetic.scala 121:25]
      end else begin
        ref_exp_diff_reg_0 <= exp_diff_out_sum_reg_1; // @[FPArithmetic.scala 128:25]
      end
    end
    if (reset) begin // @[FPArithmetic.scala 73:35]
      ref_exp_diff_reg_1 <= 8'h0; // @[FPArithmetic.scala 73:35]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_diff_reg_1 <= ref_exp_diff_reg_0; // @[FPArithmetic.scala 199:31]
    end
    if (reset) begin // @[FPArithmetic.scala 73:35]
      ref_exp_diff_reg_2 <= 8'h0; // @[FPArithmetic.scala 73:35]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_diff_reg_2 <= ref_exp_diff_reg_1; // @[FPArithmetic.scala 199:31]
    end
    if (reset) begin // @[FPArithmetic.scala 73:35]
      ref_exp_diff_reg_3 <= 8'h0; // @[FPArithmetic.scala 73:35]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_diff_reg_3 <= ref_exp_diff_reg_2; // @[FPArithmetic.scala 199:31]
    end
    if (reset) begin // @[FPArithmetic.scala 73:35]
      ref_exp_diff_reg_4 <= 8'h0; // @[FPArithmetic.scala 73:35]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_diff_reg_4 <= ref_exp_diff_reg_3; // @[FPArithmetic.scala 199:31]
    end
    if (reset) begin // @[FPArithmetic.scala 73:35]
      ref_exp_diff_reg_5 <= 8'h0; // @[FPArithmetic.scala 73:35]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_diff_reg_5 <= ref_exp_diff_reg_4; // @[FPArithmetic.scala 199:31]
    end
    if (reset) begin // @[FPArithmetic.scala 73:35]
      ref_exp_diff_reg_6 <= 8'h0; // @[FPArithmetic.scala 73:35]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_diff_reg_6 <= ref_exp_diff_reg_5; // @[FPArithmetic.scala 199:31]
    end
    if (reset) begin // @[FPArithmetic.scala 73:35]
      ref_exp_diff_reg_7 <= 8'h0; // @[FPArithmetic.scala 73:35]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_exp_diff_reg_7 <= ref_exp_diff_reg_6; // @[FPArithmetic.scala 199:31]
    end
    if (reset) begin // @[FPArithmetic.scala 75:41]
      frac_adder_out_sum_reg_0 <= 24'h0; // @[FPArithmetic.scala 75:41]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      frac_adder_out_sum_reg_0 <= frac_adder_io_out_s; // @[FPArithmetic.scala 183:33]
    end
    if (reset) begin // @[FPArithmetic.scala 75:41]
      frac_adder_out_sum_reg_1 <= 24'h0; // @[FPArithmetic.scala 75:41]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      frac_adder_out_sum_reg_1 <= frac_adder_out_sum_reg_0; // @[FPArithmetic.scala 208:37]
    end
    if (reset) begin // @[FPArithmetic.scala 75:41]
      frac_adder_out_sum_reg_2 <= 24'h0; // @[FPArithmetic.scala 75:41]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      frac_adder_out_sum_reg_2 <= frac_adder_out_sum_reg_1; // @[FPArithmetic.scala 208:37]
    end
    if (reset) begin // @[FPArithmetic.scala 76:43]
      frac_adder_out_carry_reg_0 <= 1'h0; // @[FPArithmetic.scala 76:43]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      frac_adder_out_carry_reg_0 <= frac_adder_io_out_c; // @[FPArithmetic.scala 184:35]
    end
    if (reset) begin // @[FPArithmetic.scala 82:31]
      new_sign_reg_0 <= 1'h0; // @[FPArithmetic.scala 82:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      new_sign_reg_0 <= new_sign_wire; // @[FPArithmetic.scala 180:23]
    end
    if (reset) begin // @[FPArithmetic.scala 82:31]
      new_sign_reg_1 <= 1'h0; // @[FPArithmetic.scala 82:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      new_sign_reg_1 <= new_sign_reg_0; // @[FPArithmetic.scala 204:27]
    end
    if (reset) begin // @[FPArithmetic.scala 82:31]
      new_sign_reg_2 <= 1'h0; // @[FPArithmetic.scala 82:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      new_sign_reg_2 <= new_sign_reg_1; // @[FPArithmetic.scala 204:27]
    end
    if (reset) begin // @[FPArithmetic.scala 82:31]
      new_sign_reg_3 <= 1'h0; // @[FPArithmetic.scala 82:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      new_sign_reg_3 <= new_sign_reg_2; // @[FPArithmetic.scala 204:27]
    end
    if (reset) begin // @[FPArithmetic.scala 82:31]
      new_sign_reg_4 <= 1'h0; // @[FPArithmetic.scala 82:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      new_sign_reg_4 <= new_sign_reg_3; // @[FPArithmetic.scala 204:27]
    end
    if (reset) begin // @[FPArithmetic.scala 82:31]
      new_sign_reg_5 <= 1'h0; // @[FPArithmetic.scala 82:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 223:20]
      if (input_a_reg_10[30:0] == 31'h0 & input_b_reg_10[30:0] == 31'h0) begin // @[FPArithmetic.scala 224:86]
        new_sign_reg_5 <= 1'h0; // @[FPArithmetic.scala 225:25]
      end else if (ref_exp_diff_reg_7 >= 8'h17) begin // @[FPArithmetic.scala 228:53]
        new_sign_reg_5 <= ref_sign_reg_7; // @[FPArithmetic.scala 229:25]
      end else begin
        new_sign_reg_5 <= _GEN_154;
      end
    end
    new_frac_reg_0 <= _GEN_170[22:0]; // @[FPArithmetic.scala 83:{31,31}]
    new_exp_reg_0 <= _GEN_171[7:0]; // @[FPArithmetic.scala 84:{30,30}]
    if (reset) begin // @[FPArithmetic.scala 89:36]
      noPostProcess_reg_0 <= 1'h0; // @[FPArithmetic.scala 89:36]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      noPostProcess_reg_0 <= noPostProcess_wire; // @[FPArithmetic.scala 181:28]
    end
    if (reset) begin // @[FPArithmetic.scala 89:36]
      noPostProcess_reg_1 <= 1'h0; // @[FPArithmetic.scala 89:36]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      noPostProcess_reg_1 <= noPostProcess_reg_0; // @[FPArithmetic.scala 202:32]
    end
    if (reset) begin // @[FPArithmetic.scala 89:36]
      noPostProcess_reg_2 <= 1'h0; // @[FPArithmetic.scala 89:36]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      noPostProcess_reg_2 <= noPostProcess_reg_1; // @[FPArithmetic.scala 202:32]
    end
    if (reset) begin // @[FPArithmetic.scala 89:36]
      noPostProcess_reg_3 <= 1'h0; // @[FPArithmetic.scala 89:36]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      noPostProcess_reg_3 <= noPostProcess_reg_2; // @[FPArithmetic.scala 202:32]
    end
    if (reset) begin // @[FPArithmetic.scala 89:36]
      noPostProcess_reg_4 <= 1'h0; // @[FPArithmetic.scala 89:36]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      noPostProcess_reg_4 <= noPostProcess_reg_3; // @[FPArithmetic.scala 202:32]
    end
    if (reset) begin // @[FPArithmetic.scala 90:45]
      postProcessInstruction_reg_0 <= 1'h0; // @[FPArithmetic.scala 90:45]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      postProcessInstruction_reg_0 <= postProcessInstruction_wire; // @[FPArithmetic.scala 182:37]
    end
    if (reset) begin // @[FPArithmetic.scala 90:45]
      postProcessInstruction_reg_1 <= 1'h0; // @[FPArithmetic.scala 90:45]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      postProcessInstruction_reg_1 <= postProcessInstruction_reg_0; // @[FPArithmetic.scala 203:41]
    end
    if (reset) begin // @[FPArithmetic.scala 90:45]
      postProcessInstruction_reg_2 <= 1'h0; // @[FPArithmetic.scala 90:45]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      postProcessInstruction_reg_2 <= postProcessInstruction_reg_1; // @[FPArithmetic.scala 203:41]
    end
    if (reset) begin // @[FPArithmetic.scala 90:45]
      postProcessInstruction_reg_3 <= 1'h0; // @[FPArithmetic.scala 90:45]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      postProcessInstruction_reg_3 <= postProcessInstruction_reg_2; // @[FPArithmetic.scala 203:41]
    end
    if (reset) begin // @[FPArithmetic.scala 90:45]
      postProcessInstruction_reg_4 <= 1'h0; // @[FPArithmetic.scala 90:45]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      postProcessInstruction_reg_4 <= postProcessInstruction_reg_3; // @[FPArithmetic.scala 203:41]
    end
    if (reset) begin // @[FPArithmetic.scala 92:41]
      ref_frac_adder_sum_reg_0 <= 24'h0; // @[FPArithmetic.scala 92:41]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      if (new_sign_reg_1 & ^_ref_frac_adder_sum_wire_T) begin // @[FPArithmetic.scala 157:35]
        ref_frac_adder_sum_reg_0 <= cmpl_frac_adder_out_sum_reg_0;
      end else begin
        ref_frac_adder_sum_reg_0 <= frac_adder_out_sum_reg_2;
      end
    end
    if (reset) begin // @[FPArithmetic.scala 92:41]
      ref_frac_adder_sum_reg_1 <= 24'h0; // @[FPArithmetic.scala 92:41]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_frac_adder_sum_reg_1 <= ref_frac_adder_sum_reg_0; // @[FPArithmetic.scala 207:37]
    end
    if (reset) begin // @[FPArithmetic.scala 92:41]
      ref_frac_adder_sum_reg_2 <= 24'h0; // @[FPArithmetic.scala 92:41]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      ref_frac_adder_sum_reg_2 <= ref_frac_adder_sum_reg_1; // @[FPArithmetic.scala 207:37]
    end
    if (reset) begin // @[FPArithmetic.scala 94:33]
      leadingOne_reg_0 <= 6'h0; // @[FPArithmetic.scala 94:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      leadingOne_reg_0 <= leadingOne_wire; // @[FPArithmetic.scala 186:25]
    end
    if (reset) begin // @[FPArithmetic.scala 94:33]
      leadingOne_reg_1 <= 6'h0; // @[FPArithmetic.scala 94:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      leadingOne_reg_1 <= leadingOne_reg_0; // @[FPArithmetic.scala 216:29]
    end
    if (reset) begin // @[FPArithmetic.scala 96:30]
      input_a_reg_0 <= 32'h0; // @[FPArithmetic.scala 96:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_a_reg_0 <= io_in_a; // @[FPArithmetic.scala 167:22]
    end
    if (reset) begin // @[FPArithmetic.scala 96:30]
      input_a_reg_1 <= 32'h0; // @[FPArithmetic.scala 96:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_a_reg_1 <= input_a_reg_0; // @[FPArithmetic.scala 192:26]
    end
    if (reset) begin // @[FPArithmetic.scala 96:30]
      input_a_reg_2 <= 32'h0; // @[FPArithmetic.scala 96:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_a_reg_2 <= input_a_reg_1; // @[FPArithmetic.scala 192:26]
    end
    if (reset) begin // @[FPArithmetic.scala 96:30]
      input_a_reg_3 <= 32'h0; // @[FPArithmetic.scala 96:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_a_reg_3 <= input_a_reg_2; // @[FPArithmetic.scala 192:26]
    end
    if (reset) begin // @[FPArithmetic.scala 96:30]
      input_a_reg_4 <= 32'h0; // @[FPArithmetic.scala 96:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_a_reg_4 <= input_a_reg_3; // @[FPArithmetic.scala 192:26]
    end
    if (reset) begin // @[FPArithmetic.scala 96:30]
      input_a_reg_5 <= 32'h0; // @[FPArithmetic.scala 96:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_a_reg_5 <= input_a_reg_4; // @[FPArithmetic.scala 192:26]
    end
    if (reset) begin // @[FPArithmetic.scala 96:30]
      input_a_reg_6 <= 32'h0; // @[FPArithmetic.scala 96:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_a_reg_6 <= input_a_reg_5; // @[FPArithmetic.scala 192:26]
    end
    if (reset) begin // @[FPArithmetic.scala 96:30]
      input_a_reg_7 <= 32'h0; // @[FPArithmetic.scala 96:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_a_reg_7 <= input_a_reg_6; // @[FPArithmetic.scala 192:26]
    end
    if (reset) begin // @[FPArithmetic.scala 96:30]
      input_a_reg_8 <= 32'h0; // @[FPArithmetic.scala 96:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_a_reg_8 <= input_a_reg_7; // @[FPArithmetic.scala 192:26]
    end
    if (reset) begin // @[FPArithmetic.scala 96:30]
      input_a_reg_9 <= 32'h0; // @[FPArithmetic.scala 96:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_a_reg_9 <= input_a_reg_8; // @[FPArithmetic.scala 192:26]
    end
    if (reset) begin // @[FPArithmetic.scala 96:30]
      input_a_reg_10 <= 32'h0; // @[FPArithmetic.scala 96:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_a_reg_10 <= input_a_reg_9; // @[FPArithmetic.scala 192:26]
    end
    if (reset) begin // @[FPArithmetic.scala 97:30]
      input_b_reg_0 <= 32'h0; // @[FPArithmetic.scala 97:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_b_reg_0 <= io_in_b; // @[FPArithmetic.scala 168:22]
    end
    if (reset) begin // @[FPArithmetic.scala 97:30]
      input_b_reg_1 <= 32'h0; // @[FPArithmetic.scala 97:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_b_reg_1 <= input_b_reg_0; // @[FPArithmetic.scala 193:26]
    end
    if (reset) begin // @[FPArithmetic.scala 97:30]
      input_b_reg_2 <= 32'h0; // @[FPArithmetic.scala 97:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_b_reg_2 <= input_b_reg_1; // @[FPArithmetic.scala 193:26]
    end
    if (reset) begin // @[FPArithmetic.scala 97:30]
      input_b_reg_3 <= 32'h0; // @[FPArithmetic.scala 97:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_b_reg_3 <= input_b_reg_2; // @[FPArithmetic.scala 193:26]
    end
    if (reset) begin // @[FPArithmetic.scala 97:30]
      input_b_reg_4 <= 32'h0; // @[FPArithmetic.scala 97:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_b_reg_4 <= input_b_reg_3; // @[FPArithmetic.scala 193:26]
    end
    if (reset) begin // @[FPArithmetic.scala 97:30]
      input_b_reg_5 <= 32'h0; // @[FPArithmetic.scala 97:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_b_reg_5 <= input_b_reg_4; // @[FPArithmetic.scala 193:26]
    end
    if (reset) begin // @[FPArithmetic.scala 97:30]
      input_b_reg_6 <= 32'h0; // @[FPArithmetic.scala 97:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_b_reg_6 <= input_b_reg_5; // @[FPArithmetic.scala 193:26]
    end
    if (reset) begin // @[FPArithmetic.scala 97:30]
      input_b_reg_7 <= 32'h0; // @[FPArithmetic.scala 97:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_b_reg_7 <= input_b_reg_6; // @[FPArithmetic.scala 193:26]
    end
    if (reset) begin // @[FPArithmetic.scala 97:30]
      input_b_reg_8 <= 32'h0; // @[FPArithmetic.scala 97:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_b_reg_8 <= input_b_reg_7; // @[FPArithmetic.scala 193:26]
    end
    if (reset) begin // @[FPArithmetic.scala 97:30]
      input_b_reg_9 <= 32'h0; // @[FPArithmetic.scala 97:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_b_reg_9 <= input_b_reg_8; // @[FPArithmetic.scala 193:26]
    end
    if (reset) begin // @[FPArithmetic.scala 97:30]
      input_b_reg_10 <= 32'h0; // @[FPArithmetic.scala 97:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      input_b_reg_10 <= input_b_reg_9; // @[FPArithmetic.scala 193:26]
    end
    if (reset) begin // @[FPArithmetic.scala 99:51]
      postProcess_exp_diff_out_sum_reg_0 <= 8'h0; // @[FPArithmetic.scala 99:51]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      postProcess_exp_diff_out_sum_reg_0 <= postProcess_exp_diff_subtractor_io_out_s; // @[FPArithmetic.scala 187:43]
    end
    if (reset) begin // @[FPArithmetic.scala 100:53]
      postProcess_exp_diff_out_carry_reg_0 <= 1'h0; // @[FPArithmetic.scala 100:53]
    end else if (io_in_en) begin // @[FPArithmetic.scala 166:19]
      postProcess_exp_diff_out_carry_reg_0 <= postProcess_exp_diff_subtractor_io_out_c; // @[FPArithmetic.scala 188:45]
    end
    if (reset) begin // @[FPArithmetic.scala 114:40]
      cmpl_subber_out_s_reg_0 <= 8'h0; // @[FPArithmetic.scala 114:40]
    end else if (io_in_en) begin // @[FPArithmetic.scala 115:19]
      cmpl_subber_out_s_reg_0 <= _cmpl_subber_out_s_reg_0_T_2; // @[FPArithmetic.scala 116:32]
    end
    if (reset) begin // @[FPArithmetic.scala 135:42]
      cmpl_frac_adder_inp_reg_0_0 <= 24'h0; // @[FPArithmetic.scala 135:42]
    end else if (io_in_en) begin // @[FPArithmetic.scala 136:19]
      cmpl_frac_adder_inp_reg_0_0 <= _cmpl_frac_adder_inp_reg_0_0_T_2; // @[FPArithmetic.scala 137:37]
    end
    if (reset) begin // @[FPArithmetic.scala 135:42]
      cmpl_frac_adder_inp_reg_0_1 <= 24'h0; // @[FPArithmetic.scala 135:42]
    end else if (io_in_en) begin // @[FPArithmetic.scala 136:19]
      cmpl_frac_adder_inp_reg_0_1 <= _cmpl_frac_adder_inp_reg_0_1_T_2; // @[FPArithmetic.scala 138:37]
    end
    if (reset) begin // @[FPArithmetic.scala 151:46]
      cmpl_frac_adder_out_sum_reg_0 <= 24'h0; // @[FPArithmetic.scala 151:46]
    end else if (io_in_en) begin // @[FPArithmetic.scala 152:19]
      cmpl_frac_adder_out_sum_reg_0 <= _cmpl_frac_adder_out_sum_reg_0_T_2; // @[FPArithmetic.scala 153:38]
    end
    if (reset) begin // @[FPArithmetic.scala 221:33]
      output_sum_reg <= 32'h0; // @[FPArithmetic.scala 221:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 223:20]
      output_sum_reg <= _output_sum_reg_T_1; // @[FPArithmetic.scala 260:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sign_reg_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sign_reg_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sign_reg_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  sign_reg_1_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  sign_reg_2_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  sign_reg_2_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  sign_reg_3_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sign_reg_3_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sign_reg_4_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sign_reg_4_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  sign_reg_5_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  sign_reg_5_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  sign_reg_6_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  sign_reg_6_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  sign_reg_7_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  sign_reg_7_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  sign_reg_8_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  sign_reg_8_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  sign_reg_9_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sign_reg_9_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  sign_reg_10_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  sign_reg_10_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  exp_reg_0_0 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  exp_reg_0_1 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  exp_reg_1_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  exp_reg_1_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  exp_reg_2_0 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  exp_reg_2_1 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  frac_reg_0_0 = _RAND_28[22:0];
  _RAND_29 = {1{`RANDOM}};
  frac_reg_0_1 = _RAND_29[22:0];
  _RAND_30 = {1{`RANDOM}};
  frac_reg_1_0 = _RAND_30[22:0];
  _RAND_31 = {1{`RANDOM}};
  frac_reg_1_1 = _RAND_31[22:0];
  _RAND_32 = {1{`RANDOM}};
  frac_reg_2_0 = _RAND_32[22:0];
  _RAND_33 = {1{`RANDOM}};
  frac_reg_2_1 = _RAND_33[22:0];
  _RAND_34 = {1{`RANDOM}};
  whole_frac_reg_0_0 = _RAND_34[23:0];
  _RAND_35 = {1{`RANDOM}};
  whole_frac_reg_0_1 = _RAND_35[23:0];
  _RAND_36 = {1{`RANDOM}};
  whole_frac_reg_1_0 = _RAND_36[23:0];
  _RAND_37 = {1{`RANDOM}};
  whole_frac_reg_1_1 = _RAND_37[23:0];
  _RAND_38 = {1{`RANDOM}};
  whole_frac_reg_2_0 = _RAND_38[23:0];
  _RAND_39 = {1{`RANDOM}};
  whole_frac_reg_2_1 = _RAND_39[23:0];
  _RAND_40 = {1{`RANDOM}};
  exp_diff_out_sum_reg_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  exp_diff_out_sum_reg_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  exp_diff_out_carry_reg_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  exp_diff_out_carry_reg_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  frac_adder_inp_reg_0_0 = _RAND_44[23:0];
  _RAND_45 = {1{`RANDOM}};
  frac_adder_inp_reg_0_1 = _RAND_45[23:0];
  _RAND_46 = {1{`RANDOM}};
  frac_adder_inp_reg_1_0 = _RAND_46[23:0];
  _RAND_47 = {1{`RANDOM}};
  frac_adder_inp_reg_1_1 = _RAND_47[23:0];
  _RAND_48 = {1{`RANDOM}};
  ref_sign_reg_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  ref_sign_reg_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  ref_sign_reg_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  ref_sign_reg_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  ref_sign_reg_4 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  ref_sign_reg_5 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  ref_sign_reg_6 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  ref_sign_reg_7 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  ref_frac_reg_0 = _RAND_56[22:0];
  _RAND_57 = {1{`RANDOM}};
  ref_frac_reg_1 = _RAND_57[22:0];
  _RAND_58 = {1{`RANDOM}};
  ref_frac_reg_2 = _RAND_58[22:0];
  _RAND_59 = {1{`RANDOM}};
  ref_frac_reg_3 = _RAND_59[22:0];
  _RAND_60 = {1{`RANDOM}};
  ref_frac_reg_4 = _RAND_60[22:0];
  _RAND_61 = {1{`RANDOM}};
  ref_frac_reg_5 = _RAND_61[22:0];
  _RAND_62 = {1{`RANDOM}};
  ref_frac_reg_6 = _RAND_62[22:0];
  _RAND_63 = {1{`RANDOM}};
  ref_frac_reg_7 = _RAND_63[22:0];
  _RAND_64 = {1{`RANDOM}};
  ref_exp_reg_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  ref_exp_reg_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  ref_exp_reg_2 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  ref_exp_reg_3 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  ref_exp_reg_4 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  ref_exp_reg_5 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  ref_exp_reg_6 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  ref_exp_reg_7 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  ref_exp_diff_reg_0 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  ref_exp_diff_reg_1 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  ref_exp_diff_reg_2 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  ref_exp_diff_reg_3 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  ref_exp_diff_reg_4 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  ref_exp_diff_reg_5 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  ref_exp_diff_reg_6 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  ref_exp_diff_reg_7 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  frac_adder_out_sum_reg_0 = _RAND_80[23:0];
  _RAND_81 = {1{`RANDOM}};
  frac_adder_out_sum_reg_1 = _RAND_81[23:0];
  _RAND_82 = {1{`RANDOM}};
  frac_adder_out_sum_reg_2 = _RAND_82[23:0];
  _RAND_83 = {1{`RANDOM}};
  frac_adder_out_carry_reg_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  new_sign_reg_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  new_sign_reg_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  new_sign_reg_2 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  new_sign_reg_3 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  new_sign_reg_4 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  new_sign_reg_5 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  new_frac_reg_0 = _RAND_90[22:0];
  _RAND_91 = {1{`RANDOM}};
  new_exp_reg_0 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  noPostProcess_reg_0 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  noPostProcess_reg_1 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  noPostProcess_reg_2 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  noPostProcess_reg_3 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  noPostProcess_reg_4 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  postProcessInstruction_reg_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  postProcessInstruction_reg_1 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  postProcessInstruction_reg_2 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  postProcessInstruction_reg_3 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  postProcessInstruction_reg_4 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  ref_frac_adder_sum_reg_0 = _RAND_102[23:0];
  _RAND_103 = {1{`RANDOM}};
  ref_frac_adder_sum_reg_1 = _RAND_103[23:0];
  _RAND_104 = {1{`RANDOM}};
  ref_frac_adder_sum_reg_2 = _RAND_104[23:0];
  _RAND_105 = {1{`RANDOM}};
  leadingOne_reg_0 = _RAND_105[5:0];
  _RAND_106 = {1{`RANDOM}};
  leadingOne_reg_1 = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  input_a_reg_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  input_a_reg_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  input_a_reg_2 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  input_a_reg_3 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  input_a_reg_4 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  input_a_reg_5 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  input_a_reg_6 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  input_a_reg_7 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  input_a_reg_8 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  input_a_reg_9 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  input_a_reg_10 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  input_b_reg_0 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  input_b_reg_1 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  input_b_reg_2 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  input_b_reg_3 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  input_b_reg_4 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  input_b_reg_5 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  input_b_reg_6 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  input_b_reg_7 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  input_b_reg_8 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  input_b_reg_9 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  input_b_reg_10 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  postProcess_exp_diff_out_sum_reg_0 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  postProcess_exp_diff_out_carry_reg_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  cmpl_subber_out_s_reg_0 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  cmpl_frac_adder_inp_reg_0_0 = _RAND_132[23:0];
  _RAND_133 = {1{`RANDOM}};
  cmpl_frac_adder_inp_reg_0_1 = _RAND_133[23:0];
  _RAND_134 = {1{`RANDOM}};
  cmpl_frac_adder_out_sum_reg_0 = _RAND_134[23:0];
  _RAND_135 = {1{`RANDOM}};
  output_sum_reg = _RAND_135[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexAdder_bw32(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input         io_in_valid,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im,
  output        io_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  FP_adder_bw32_clock; // @[FPComplex.scala 27:42]
  wire  FP_adder_bw32_reset; // @[FPComplex.scala 27:42]
  wire  FP_adder_bw32_io_in_en; // @[FPComplex.scala 27:42]
  wire [31:0] FP_adder_bw32_io_in_a; // @[FPComplex.scala 27:42]
  wire [31:0] FP_adder_bw32_io_in_b; // @[FPComplex.scala 27:42]
  wire [31:0] FP_adder_bw32_io_out_s; // @[FPComplex.scala 27:42]
  wire  FP_adder_bw32_1_clock; // @[FPComplex.scala 27:42]
  wire  FP_adder_bw32_1_reset; // @[FPComplex.scala 27:42]
  wire  FP_adder_bw32_1_io_in_en; // @[FPComplex.scala 27:42]
  wire [31:0] FP_adder_bw32_1_io_in_a; // @[FPComplex.scala 27:42]
  wire [31:0] FP_adder_bw32_1_io_in_b; // @[FPComplex.scala 27:42]
  wire [31:0] FP_adder_bw32_1_io_out_s; // @[FPComplex.scala 27:42]
  reg  io_out_valid_r; // @[Reg.scala 16:16]
  reg  io_out_valid_r_1; // @[Reg.scala 16:16]
  reg  io_out_valid_r_2; // @[Reg.scala 16:16]
  reg  io_out_valid_r_3; // @[Reg.scala 16:16]
  reg  io_out_valid_r_4; // @[Reg.scala 16:16]
  reg  io_out_valid_r_5; // @[Reg.scala 16:16]
  reg  io_out_valid_r_6; // @[Reg.scala 16:16]
  reg  io_out_valid_r_7; // @[Reg.scala 16:16]
  reg  io_out_valid_r_8; // @[Reg.scala 16:16]
  reg  io_out_valid_r_9; // @[Reg.scala 16:16]
  reg  io_out_valid_r_10; // @[Reg.scala 16:16]
  reg  io_out_valid_r_11; // @[Reg.scala 16:16]
  reg  io_out_valid_r_12; // @[Reg.scala 16:16]
  FP_adder_bw32 FP_adder_bw32 ( // @[FPComplex.scala 27:42]
    .clock(FP_adder_bw32_clock),
    .reset(FP_adder_bw32_reset),
    .io_in_en(FP_adder_bw32_io_in_en),
    .io_in_a(FP_adder_bw32_io_in_a),
    .io_in_b(FP_adder_bw32_io_in_b),
    .io_out_s(FP_adder_bw32_io_out_s)
  );
  FP_adder_bw32 FP_adder_bw32_1 ( // @[FPComplex.scala 27:42]
    .clock(FP_adder_bw32_1_clock),
    .reset(FP_adder_bw32_1_reset),
    .io_in_en(FP_adder_bw32_1_io_in_en),
    .io_in_a(FP_adder_bw32_1_io_in_a),
    .io_in_b(FP_adder_bw32_1_io_in_b),
    .io_out_s(FP_adder_bw32_1_io_out_s)
  );
  assign io_out_s_Re = FP_adder_bw32_io_out_s; // @[FPComplex.scala 34:17]
  assign io_out_s_Im = FP_adder_bw32_1_io_out_s; // @[FPComplex.scala 35:17]
  assign io_out_valid = io_out_valid_r_12; // @[FPComplex.scala 36:18]
  assign FP_adder_bw32_clock = clock;
  assign FP_adder_bw32_reset = reset;
  assign FP_adder_bw32_io_in_en = io_in_en; // @[FPComplex.scala 28:24]
  assign FP_adder_bw32_io_in_a = io_in_a_Re; // @[FPComplex.scala 30:23]
  assign FP_adder_bw32_io_in_b = io_in_b_Re; // @[FPComplex.scala 31:23]
  assign FP_adder_bw32_1_clock = clock;
  assign FP_adder_bw32_1_reset = reset;
  assign FP_adder_bw32_1_io_in_en = io_in_en; // @[FPComplex.scala 29:24]
  assign FP_adder_bw32_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 32:23]
  assign FP_adder_bw32_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 33:23]
  always @(posedge clock) begin
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r <= io_in_valid; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_1 <= io_out_valid_r; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_2 <= io_out_valid_r_1; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_3 <= io_out_valid_r_2; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_4 <= io_out_valid_r_3; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_5 <= io_out_valid_r_4; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_6 <= io_out_valid_r_5; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_7 <= io_out_valid_r_6; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_8 <= io_out_valid_r_7; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_9 <= io_out_valid_r_8; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_10 <= io_out_valid_r_9; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_11 <= io_out_valid_r_10; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_12 <= io_out_valid_r_11; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_valid_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_out_valid_r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_out_valid_r_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  io_out_valid_r_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_out_valid_r_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  io_out_valid_r_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  io_out_valid_r_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_out_valid_r_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_out_valid_r_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  io_out_valid_r_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_out_valid_r_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  io_out_valid_r_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  io_out_valid_r_12 = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FP_subtractor_bw32(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire  FP_adder_clock; // @[FPArithmetic.scala 274:26]
  wire  FP_adder_reset; // @[FPArithmetic.scala 274:26]
  wire  FP_adder_io_in_en; // @[FPArithmetic.scala 274:26]
  wire [31:0] FP_adder_io_in_a; // @[FPArithmetic.scala 274:26]
  wire [31:0] FP_adder_io_in_b; // @[FPArithmetic.scala 274:26]
  wire [31:0] FP_adder_io_out_s; // @[FPArithmetic.scala 274:26]
  wire  _adjusted_in_b_T_1 = ~io_in_b[31]; // @[FPArithmetic.scala 276:23]
  FP_adder_bw32 FP_adder ( // @[FPArithmetic.scala 274:26]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_en(FP_adder_io_in_en),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  assign io_out_s = FP_adder_io_out_s; // @[FPArithmetic.scala 280:14]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_en = io_in_en; // @[FPArithmetic.scala 277:23]
  assign FP_adder_io_in_a = io_in_a; // @[FPArithmetic.scala 278:22]
  assign FP_adder_io_in_b = {_adjusted_in_b_T_1,io_in_b[30:0]}; // @[FPArithmetic.scala 276:41]
endmodule
module FPComplexSubtractor_bw32(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire  FP_subtractor_bw32_clock; // @[FPComplex.scala 87:47]
  wire  FP_subtractor_bw32_reset; // @[FPComplex.scala 87:47]
  wire  FP_subtractor_bw32_io_in_en; // @[FPComplex.scala 87:47]
  wire [31:0] FP_subtractor_bw32_io_in_a; // @[FPComplex.scala 87:47]
  wire [31:0] FP_subtractor_bw32_io_in_b; // @[FPComplex.scala 87:47]
  wire [31:0] FP_subtractor_bw32_io_out_s; // @[FPComplex.scala 87:47]
  wire  FP_subtractor_bw32_1_clock; // @[FPComplex.scala 87:47]
  wire  FP_subtractor_bw32_1_reset; // @[FPComplex.scala 87:47]
  wire  FP_subtractor_bw32_1_io_in_en; // @[FPComplex.scala 87:47]
  wire [31:0] FP_subtractor_bw32_1_io_in_a; // @[FPComplex.scala 87:47]
  wire [31:0] FP_subtractor_bw32_1_io_in_b; // @[FPComplex.scala 87:47]
  wire [31:0] FP_subtractor_bw32_1_io_out_s; // @[FPComplex.scala 87:47]
  FP_subtractor_bw32 FP_subtractor_bw32 ( // @[FPComplex.scala 87:47]
    .clock(FP_subtractor_bw32_clock),
    .reset(FP_subtractor_bw32_reset),
    .io_in_en(FP_subtractor_bw32_io_in_en),
    .io_in_a(FP_subtractor_bw32_io_in_a),
    .io_in_b(FP_subtractor_bw32_io_in_b),
    .io_out_s(FP_subtractor_bw32_io_out_s)
  );
  FP_subtractor_bw32 FP_subtractor_bw32_1 ( // @[FPComplex.scala 87:47]
    .clock(FP_subtractor_bw32_1_clock),
    .reset(FP_subtractor_bw32_1_reset),
    .io_in_en(FP_subtractor_bw32_1_io_in_en),
    .io_in_a(FP_subtractor_bw32_1_io_in_a),
    .io_in_b(FP_subtractor_bw32_1_io_in_b),
    .io_out_s(FP_subtractor_bw32_1_io_out_s)
  );
  assign io_out_s_Re = FP_subtractor_bw32_io_out_s; // @[FPComplex.scala 94:17]
  assign io_out_s_Im = FP_subtractor_bw32_1_io_out_s; // @[FPComplex.scala 95:17]
  assign FP_subtractor_bw32_clock = clock;
  assign FP_subtractor_bw32_reset = reset;
  assign FP_subtractor_bw32_io_in_en = io_in_en; // @[FPComplex.scala 88:29]
  assign FP_subtractor_bw32_io_in_a = io_in_a_Re; // @[FPComplex.scala 90:28]
  assign FP_subtractor_bw32_io_in_b = io_in_b_Re; // @[FPComplex.scala 91:28]
  assign FP_subtractor_bw32_1_clock = clock;
  assign FP_subtractor_bw32_1_reset = reset;
  assign FP_subtractor_bw32_1_io_in_en = io_in_en; // @[FPComplex.scala 89:29]
  assign FP_subtractor_bw32_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 92:28]
  assign FP_subtractor_bw32_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 93:28]
endmodule
module DFT_2_bw32(
  input         clock,
  input         reset,
  input         io_in_en,
  input         io_in_valid,
  input  [31:0] io_in_data_0_Re,
  input  [31:0] io_in_data_0_Im,
  input  [31:0] io_in_data_1_Re,
  input  [31:0] io_in_data_1_Im,
  output        io_out_valid,
  output [31:0] io_out_data_0_Re,
  output [31:0] io_out_data_0_Im,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  FPComplexAdder_bw32_clock; // @[DFTDesigns.scala 26:23]
  wire  FPComplexAdder_bw32_reset; // @[DFTDesigns.scala 26:23]
  wire  FPComplexAdder_bw32_io_in_en; // @[DFTDesigns.scala 26:23]
  wire [31:0] FPComplexAdder_bw32_io_in_a_Re; // @[DFTDesigns.scala 26:23]
  wire [31:0] FPComplexAdder_bw32_io_in_a_Im; // @[DFTDesigns.scala 26:23]
  wire  FPComplexAdder_bw32_io_in_valid; // @[DFTDesigns.scala 26:23]
  wire [31:0] FPComplexAdder_bw32_io_in_b_Re; // @[DFTDesigns.scala 26:23]
  wire [31:0] FPComplexAdder_bw32_io_in_b_Im; // @[DFTDesigns.scala 26:23]
  wire [31:0] FPComplexAdder_bw32_io_out_s_Re; // @[DFTDesigns.scala 26:23]
  wire [31:0] FPComplexAdder_bw32_io_out_s_Im; // @[DFTDesigns.scala 26:23]
  wire  FPComplexAdder_bw32_io_out_valid; // @[DFTDesigns.scala 26:23]
  wire  FPComplexSubtractor_bw32_clock; // @[DFTDesigns.scala 27:28]
  wire  FPComplexSubtractor_bw32_reset; // @[DFTDesigns.scala 27:28]
  wire  FPComplexSubtractor_bw32_io_in_en; // @[DFTDesigns.scala 27:28]
  wire [31:0] FPComplexSubtractor_bw32_io_in_a_Re; // @[DFTDesigns.scala 27:28]
  wire [31:0] FPComplexSubtractor_bw32_io_in_a_Im; // @[DFTDesigns.scala 27:28]
  wire [31:0] FPComplexSubtractor_bw32_io_in_b_Re; // @[DFTDesigns.scala 27:28]
  wire [31:0] FPComplexSubtractor_bw32_io_in_b_Im; // @[DFTDesigns.scala 27:28]
  wire [31:0] FPComplexSubtractor_bw32_io_out_s_Re; // @[DFTDesigns.scala 27:28]
  wire [31:0] FPComplexSubtractor_bw32_io_out_s_Im; // @[DFTDesigns.scala 27:28]
  reg  io_out_valid_r; // @[Reg.scala 16:16]
  reg [31:0] io_out_data_0_r_Re; // @[Reg.scala 16:16]
  reg [31:0] io_out_data_0_r_Im; // @[Reg.scala 16:16]
  reg [31:0] io_out_data_1_r_Re; // @[Reg.scala 16:16]
  reg [31:0] io_out_data_1_r_Im; // @[Reg.scala 16:16]
  FPComplexAdder_bw32 FPComplexAdder_bw32 ( // @[DFTDesigns.scala 26:23]
    .clock(FPComplexAdder_bw32_clock),
    .reset(FPComplexAdder_bw32_reset),
    .io_in_en(FPComplexAdder_bw32_io_in_en),
    .io_in_a_Re(FPComplexAdder_bw32_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_bw32_io_in_a_Im),
    .io_in_valid(FPComplexAdder_bw32_io_in_valid),
    .io_in_b_Re(FPComplexAdder_bw32_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_bw32_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_bw32_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_bw32_io_out_s_Im),
    .io_out_valid(FPComplexAdder_bw32_io_out_valid)
  );
  FPComplexSubtractor_bw32 FPComplexSubtractor_bw32 ( // @[DFTDesigns.scala 27:28]
    .clock(FPComplexSubtractor_bw32_clock),
    .reset(FPComplexSubtractor_bw32_reset),
    .io_in_en(FPComplexSubtractor_bw32_io_in_en),
    .io_in_a_Re(FPComplexSubtractor_bw32_io_in_a_Re),
    .io_in_a_Im(FPComplexSubtractor_bw32_io_in_a_Im),
    .io_in_b_Re(FPComplexSubtractor_bw32_io_in_b_Re),
    .io_in_b_Im(FPComplexSubtractor_bw32_io_in_b_Im),
    .io_out_s_Re(FPComplexSubtractor_bw32_io_out_s_Re),
    .io_out_s_Im(FPComplexSubtractor_bw32_io_out_s_Im)
  );
  assign io_out_valid = io_out_valid_r; // @[DFTDesigns.scala 30:18]
  assign io_out_data_0_Re = io_out_data_0_r_Re; // @[DFTDesigns.scala 37:20]
  assign io_out_data_0_Im = io_out_data_0_r_Im; // @[DFTDesigns.scala 37:20]
  assign io_out_data_1_Re = io_out_data_1_r_Re; // @[DFTDesigns.scala 38:20]
  assign io_out_data_1_Im = io_out_data_1_r_Im; // @[DFTDesigns.scala 38:20]
  assign FPComplexAdder_bw32_clock = clock;
  assign FPComplexAdder_bw32_reset = reset;
  assign FPComplexAdder_bw32_io_in_en = io_in_en; // @[DFTDesigns.scala 31:17]
  assign FPComplexAdder_bw32_io_in_a_Re = io_in_data_0_Re; // @[DFTDesigns.scala 33:16]
  assign FPComplexAdder_bw32_io_in_a_Im = io_in_data_0_Im; // @[DFTDesigns.scala 33:16]
  assign FPComplexAdder_bw32_io_in_valid = io_in_valid; // @[DFTDesigns.scala 28:20]
  assign FPComplexAdder_bw32_io_in_b_Re = io_in_data_1_Re; // @[DFTDesigns.scala 34:16]
  assign FPComplexAdder_bw32_io_in_b_Im = io_in_data_1_Im; // @[DFTDesigns.scala 34:16]
  assign FPComplexSubtractor_bw32_clock = clock;
  assign FPComplexSubtractor_bw32_reset = reset;
  assign FPComplexSubtractor_bw32_io_in_en = io_in_en; // @[DFTDesigns.scala 32:22]
  assign FPComplexSubtractor_bw32_io_in_a_Re = io_in_data_0_Re; // @[DFTDesigns.scala 35:21]
  assign FPComplexSubtractor_bw32_io_in_a_Im = io_in_data_0_Im; // @[DFTDesigns.scala 35:21]
  assign FPComplexSubtractor_bw32_io_in_b_Re = io_in_data_1_Re; // @[DFTDesigns.scala 36:21]
  assign FPComplexSubtractor_bw32_io_in_b_Im = io_in_data_1_Im; // @[DFTDesigns.scala 36:21]
  always @(posedge clock) begin
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r <= FPComplexAdder_bw32_io_out_valid; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_data_0_r_Re <= FPComplexAdder_bw32_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_data_0_r_Im <= FPComplexAdder_bw32_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_data_1_r_Re <= FPComplexSubtractor_bw32_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_data_1_r_Im <= FPComplexSubtractor_bw32_io_out_s_Im; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_valid_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_out_data_0_r_Re = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  io_out_data_0_r_Im = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_out_data_1_r_Re = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  io_out_data_1_r_Im = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DFT2_bw32(
  input         clock,
  input         reset,
  input         io_in_en,
  input         io_in_valid,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output        io_out_valid
);
  wire  DFT_2_bw32_clock; // @[DFTDesigns.scala 55:24]
  wire  DFT_2_bw32_reset; // @[DFTDesigns.scala 55:24]
  wire  DFT_2_bw32_io_in_en; // @[DFTDesigns.scala 55:24]
  wire  DFT_2_bw32_io_in_valid; // @[DFTDesigns.scala 55:24]
  wire [31:0] DFT_2_bw32_io_in_data_0_Re; // @[DFTDesigns.scala 55:24]
  wire [31:0] DFT_2_bw32_io_in_data_0_Im; // @[DFTDesigns.scala 55:24]
  wire [31:0] DFT_2_bw32_io_in_data_1_Re; // @[DFTDesigns.scala 55:24]
  wire [31:0] DFT_2_bw32_io_in_data_1_Im; // @[DFTDesigns.scala 55:24]
  wire  DFT_2_bw32_io_out_valid; // @[DFTDesigns.scala 55:24]
  wire [31:0] DFT_2_bw32_io_out_data_0_Re; // @[DFTDesigns.scala 55:24]
  wire [31:0] DFT_2_bw32_io_out_data_0_Im; // @[DFTDesigns.scala 55:24]
  wire [31:0] DFT_2_bw32_io_out_data_1_Re; // @[DFTDesigns.scala 55:24]
  wire [31:0] DFT_2_bw32_io_out_data_1_Im; // @[DFTDesigns.scala 55:24]
  DFT_2_bw32 DFT_2_bw32 ( // @[DFTDesigns.scala 55:24]
    .clock(DFT_2_bw32_clock),
    .reset(DFT_2_bw32_reset),
    .io_in_en(DFT_2_bw32_io_in_en),
    .io_in_valid(DFT_2_bw32_io_in_valid),
    .io_in_data_0_Re(DFT_2_bw32_io_in_data_0_Re),
    .io_in_data_0_Im(DFT_2_bw32_io_in_data_0_Im),
    .io_in_data_1_Re(DFT_2_bw32_io_in_data_1_Re),
    .io_in_data_1_Im(DFT_2_bw32_io_in_data_1_Im),
    .io_out_valid(DFT_2_bw32_io_out_valid),
    .io_out_data_0_Re(DFT_2_bw32_io_out_data_0_Re),
    .io_out_data_0_Im(DFT_2_bw32_io_out_data_0_Im),
    .io_out_data_1_Re(DFT_2_bw32_io_out_data_1_Re),
    .io_out_data_1_Im(DFT_2_bw32_io_out_data_1_Im)
  );
  assign io_out_0_Re = DFT_2_bw32_io_out_data_0_Re; // @[DFTDesigns.scala 59:14]
  assign io_out_0_Im = DFT_2_bw32_io_out_data_0_Im; // @[DFTDesigns.scala 59:14]
  assign io_out_1_Re = DFT_2_bw32_io_out_data_1_Re; // @[DFTDesigns.scala 59:14]
  assign io_out_1_Im = DFT_2_bw32_io_out_data_1_Im; // @[DFTDesigns.scala 59:14]
  assign io_out_valid = DFT_2_bw32_io_out_valid; // @[DFTDesigns.scala 60:20]
  assign DFT_2_bw32_clock = clock;
  assign DFT_2_bw32_reset = reset;
  assign DFT_2_bw32_io_in_en = io_in_en; // @[DFTDesigns.scala 56:18]
  assign DFT_2_bw32_io_in_valid = io_in_valid; // @[DFTDesigns.scala 57:21]
  assign DFT_2_bw32_io_in_data_0_Re = io_in_0_Re; // @[DFTDesigns.scala 58:20]
  assign DFT_2_bw32_io_in_data_0_Im = io_in_0_Im; // @[DFTDesigns.scala 58:20]
  assign DFT_2_bw32_io_in_data_1_Re = io_in_1_Re; // @[DFTDesigns.scala 58:20]
  assign DFT_2_bw32_io_in_data_1_Im = io_in_1_Im; // @[DFTDesigns.scala 58:20]
endmodule
module simple_RAM_depth2_bw64(
  input         clock,
  input         io_in_addr,
  input  [63:0] io_in_data,
  input         io_in_en,
  input         io_in_we,
  output [63:0] io_out_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] smem [0:1]; // @[PaddingDesigns.scala 42:27]
  wire  smem_io_out_data_MPORT_en; // @[PaddingDesigns.scala 42:27]
  wire  smem_io_out_data_MPORT_addr; // @[PaddingDesigns.scala 42:27]
  wire [63:0] smem_io_out_data_MPORT_data; // @[PaddingDesigns.scala 42:27]
  wire [63:0] smem_MPORT_data; // @[PaddingDesigns.scala 42:27]
  wire  smem_MPORT_addr; // @[PaddingDesigns.scala 42:27]
  wire  smem_MPORT_mask; // @[PaddingDesigns.scala 42:27]
  wire  smem_MPORT_en; // @[PaddingDesigns.scala 42:27]
  reg  smem_io_out_data_MPORT_en_pipe_0;
  reg  smem_io_out_data_MPORT_addr_pipe_0;
  wire  _io_out_data_T = ~io_in_we; // @[PaddingDesigns.scala 45:52]
  assign smem_io_out_data_MPORT_en = smem_io_out_data_MPORT_en_pipe_0;
  assign smem_io_out_data_MPORT_addr = smem_io_out_data_MPORT_addr_pipe_0;
  assign smem_io_out_data_MPORT_data = smem[smem_io_out_data_MPORT_addr]; // @[PaddingDesigns.scala 42:27]
  assign smem_MPORT_data = io_in_data;
  assign smem_MPORT_addr = io_in_addr;
  assign smem_MPORT_mask = 1'h1;
  assign smem_MPORT_en = io_in_we & io_in_en;
  assign io_out_data = smem_io_out_data_MPORT_data; // @[PaddingDesigns.scala 45:17]
  always @(posedge clock) begin
    if (smem_MPORT_en & smem_MPORT_mask) begin
      smem[smem_MPORT_addr] <= smem_MPORT_data; // @[PaddingDesigns.scala 42:27]
    end
    smem_io_out_data_MPORT_en_pipe_0 <= io_in_en & _io_out_data_T;
    if (io_in_en & _io_out_data_T) begin
      smem_io_out_data_MPORT_addr_pipe_0 <= io_in_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    smem[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  smem_io_out_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  smem_io_out_data_MPORT_addr_pipe_0 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RAM_n2_bw64(
  input         clock,
  input         io_in_en,
  input         io_in_valid,
  input  [63:0] io_in_data,
  input         io_in_we,
  input  [1:0]  io_in_addr,
  output [63:0] io_out_data
);
  wire  simple_RAM_depth2_bw64_clock; // @[PermutationDesigns.scala 276:22]
  wire  simple_RAM_depth2_bw64_io_in_addr; // @[PermutationDesigns.scala 276:22]
  wire [63:0] simple_RAM_depth2_bw64_io_in_data; // @[PermutationDesigns.scala 276:22]
  wire  simple_RAM_depth2_bw64_io_in_en; // @[PermutationDesigns.scala 276:22]
  wire  simple_RAM_depth2_bw64_io_in_we; // @[PermutationDesigns.scala 276:22]
  wire [63:0] simple_RAM_depth2_bw64_io_out_data; // @[PermutationDesigns.scala 276:22]
  wire [63:0] _GEN_0 = io_in_valid ? io_in_data : 64'h0; // @[PermutationDesigns.scala 277:18 286:27 287:24]
  wire [1:0] _GEN_2 = io_in_valid ? io_in_addr : 2'h0; // @[PermutationDesigns.scala 278:18 286:27 289:24]
  wire [63:0] _GEN_3 = io_in_we ? _GEN_0 : 64'h0; // @[PermutationDesigns.scala 277:18 285:21]
  wire  _GEN_4 = io_in_we & io_in_valid; // @[PermutationDesigns.scala 285:21 293:20]
  wire [1:0] _GEN_5 = io_in_we ? _GEN_2 : io_in_addr; // @[PermutationDesigns.scala 285:21 294:22]
  wire [1:0] _GEN_9 = io_in_en ? _GEN_5 : 2'h0; // @[PermutationDesigns.scala 278:18 284:19]
  simple_RAM_depth2_bw64 simple_RAM_depth2_bw64 ( // @[PermutationDesigns.scala 276:22]
    .clock(simple_RAM_depth2_bw64_clock),
    .io_in_addr(simple_RAM_depth2_bw64_io_in_addr),
    .io_in_data(simple_RAM_depth2_bw64_io_in_data),
    .io_in_en(simple_RAM_depth2_bw64_io_in_en),
    .io_in_we(simple_RAM_depth2_bw64_io_in_we),
    .io_out_data(simple_RAM_depth2_bw64_io_out_data)
  );
  assign io_out_data = simple_RAM_depth2_bw64_io_out_data; // @[PermutationDesigns.scala 283:17]
  assign simple_RAM_depth2_bw64_clock = clock;
  assign simple_RAM_depth2_bw64_io_in_addr = _GEN_9[0];
  assign simple_RAM_depth2_bw64_io_in_data = io_in_en ? _GEN_3 : 64'h0; // @[PermutationDesigns.scala 277:18 284:19]
  assign simple_RAM_depth2_bw64_io_in_en = io_in_en; // @[PermutationDesigns.scala 280:16]
  assign simple_RAM_depth2_bw64_io_in_we = io_in_en & _GEN_4; // @[PermutationDesigns.scala 279:16 284:19]
endmodule
module RAM_Block_N32_w16_bw64(
  input         clock,
  input  [1:0]  io_in_raddr,
  input  [1:0]  io_in_waddr,
  input  [63:0] io_in_data,
  input         io_in_offset_switch,
  input         io_in_valid,
  input         io_in_en,
  output [63:0] io_out_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_n2_bw64_clock; // @[PermutationDesigns.scala 249:35]
  wire  RAM_n2_bw64_io_in_en; // @[PermutationDesigns.scala 249:35]
  wire  RAM_n2_bw64_io_in_valid; // @[PermutationDesigns.scala 249:35]
  wire [63:0] RAM_n2_bw64_io_in_data; // @[PermutationDesigns.scala 249:35]
  wire  RAM_n2_bw64_io_in_we; // @[PermutationDesigns.scala 249:35]
  wire [1:0] RAM_n2_bw64_io_in_addr; // @[PermutationDesigns.scala 249:35]
  wire [63:0] RAM_n2_bw64_io_out_data; // @[PermutationDesigns.scala 249:35]
  wire  RAM_n2_bw64_1_clock; // @[PermutationDesigns.scala 249:35]
  wire  RAM_n2_bw64_1_io_in_en; // @[PermutationDesigns.scala 249:35]
  wire  RAM_n2_bw64_1_io_in_valid; // @[PermutationDesigns.scala 249:35]
  wire [63:0] RAM_n2_bw64_1_io_in_data; // @[PermutationDesigns.scala 249:35]
  wire  RAM_n2_bw64_1_io_in_we; // @[PermutationDesigns.scala 249:35]
  wire [1:0] RAM_n2_bw64_1_io_in_addr; // @[PermutationDesigns.scala 249:35]
  wire [63:0] RAM_n2_bw64_1_io_out_data; // @[PermutationDesigns.scala 249:35]
  reg  offset_switch_reg; // @[Reg.scala 16:16]
  wire  _T_1 = ~io_in_offset_switch; // @[PermutationDesigns.scala 258:21]
  RAM_n2_bw64 RAM_n2_bw64 ( // @[PermutationDesigns.scala 249:35]
    .clock(RAM_n2_bw64_clock),
    .io_in_en(RAM_n2_bw64_io_in_en),
    .io_in_valid(RAM_n2_bw64_io_in_valid),
    .io_in_data(RAM_n2_bw64_io_in_data),
    .io_in_we(RAM_n2_bw64_io_in_we),
    .io_in_addr(RAM_n2_bw64_io_in_addr),
    .io_out_data(RAM_n2_bw64_io_out_data)
  );
  RAM_n2_bw64 RAM_n2_bw64_1 ( // @[PermutationDesigns.scala 249:35]
    .clock(RAM_n2_bw64_1_clock),
    .io_in_en(RAM_n2_bw64_1_io_in_en),
    .io_in_valid(RAM_n2_bw64_1_io_in_valid),
    .io_in_data(RAM_n2_bw64_1_io_in_data),
    .io_in_we(RAM_n2_bw64_1_io_in_we),
    .io_in_addr(RAM_n2_bw64_1_io_in_addr),
    .io_out_data(RAM_n2_bw64_1_io_out_data)
  );
  assign io_out_data = offset_switch_reg ? RAM_n2_bw64_io_out_data : RAM_n2_bw64_1_io_out_data; // @[PermutationDesigns.scala 262:23]
  assign RAM_n2_bw64_clock = clock;
  assign RAM_n2_bw64_io_in_en = io_in_en; // @[PermutationDesigns.scala 256:18]
  assign RAM_n2_bw64_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 257:21]
  assign RAM_n2_bw64_io_in_data = io_in_data; // @[PermutationDesigns.scala 259:20]
  assign RAM_n2_bw64_io_in_we = ~io_in_offset_switch; // @[PermutationDesigns.scala 258:21]
  assign RAM_n2_bw64_io_in_addr = _T_1 ? io_in_waddr : io_in_raddr; // @[PermutationDesigns.scala 260:26]
  assign RAM_n2_bw64_1_clock = clock;
  assign RAM_n2_bw64_1_io_in_en = io_in_en; // @[PermutationDesigns.scala 251:18]
  assign RAM_n2_bw64_1_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 252:21]
  assign RAM_n2_bw64_1_io_in_data = io_in_data; // @[PermutationDesigns.scala 254:20]
  assign RAM_n2_bw64_1_io_in_we = io_in_offset_switch; // @[PermutationDesigns.scala 253:18]
  assign RAM_n2_bw64_1_io_in_addr = io_in_offset_switch ? io_in_waddr : io_in_raddr; // @[PermutationDesigns.scala 255:26]
  always @(posedge clock) begin
    if (io_in_en) begin // @[Reg.scala 17:18]
      offset_switch_reg <= io_in_offset_switch; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_switch_reg = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0(
  input   io_in_cnt,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15
);
  assign io_out_0 = io_in_cnt; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_1 = io_in_cnt ? 1'h0 : 1'h1; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_2 = io_in_cnt; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_3 = io_in_cnt ? 1'h0 : 1'h1; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_4 = io_in_cnt; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_5 = io_in_cnt ? 1'h0 : 1'h1; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_6 = io_in_cnt; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_7 = io_in_cnt ? 1'h0 : 1'h1; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_8 = io_in_cnt; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_9 = io_in_cnt ? 1'h0 : 1'h1; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_10 = io_in_cnt; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_11 = io_in_cnt ? 1'h0 : 1'h1; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_12 = io_in_cnt; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_13 = io_in_cnt ? 1'h0 : 1'h1; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_14 = io_in_cnt; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_15 = io_in_cnt ? 1'h0 : 1'h1; // @[PermutationDesigns.scala 229:{31,31}]
endmodule
module Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1(
  input        clock,
  input        io_in_en,
  input        io_in_cnt,
  output [3:0] io_out_0,
  output [3:0] io_out_1,
  output [3:0] io_out_2,
  output [3:0] io_out_3,
  output [3:0] io_out_4,
  output [3:0] io_out_5,
  output [3:0] io_out_6,
  output [3:0] io_out_7,
  output [3:0] io_out_8,
  output [3:0] io_out_9,
  output [3:0] io_out_10,
  output [3:0] io_out_11,
  output [3:0] io_out_12,
  output [3:0] io_out_13,
  output [3:0] io_out_14,
  output [3:0] io_out_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] out_reg_data_r; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_1; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_2; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_3; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_4; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_5; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_6; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_7; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_8; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_9; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_10; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_11; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_12; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_13; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_14; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_15; // @[Reg.scala 16:16]
  assign io_out_0 = out_reg_data_r; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_1 = out_reg_data_r_1; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_2 = out_reg_data_r_2; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_3 = out_reg_data_r_3; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_4 = out_reg_data_r_4; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_5 = out_reg_data_r_5; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_6 = out_reg_data_r_6; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_7 = out_reg_data_r_7; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_8 = out_reg_data_r_8; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_9 = out_reg_data_r_9; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_10 = out_reg_data_r_10; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_11 = out_reg_data_r_11; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_12 = out_reg_data_r_12; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_13 = out_reg_data_r_13; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_14 = out_reg_data_r_14; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_15 = out_reg_data_r_15; // @[PermutationDesigns.scala 229:{31,31}]
  always @(posedge clock) begin
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r <= 4'h1; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r <= 4'h0;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_1 <= 4'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_1 <= 4'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_2 <= 4'h9; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_2 <= 4'h8;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_3 <= 4'h8; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_3 <= 4'h9;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_4 <= 4'h5; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_4 <= 4'h4;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_5 <= 4'h4; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_5 <= 4'h5;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_6 <= 4'hd; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_6 <= 4'hc;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_7 <= 4'hc; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_7 <= 4'hd;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_8 <= 4'h3; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_8 <= 4'h2;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_9 <= 4'h2; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_9 <= 4'h3;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_10 <= 4'hb; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_10 <= 4'ha;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_11 <= 4'ha; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_11 <= 4'hb;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_12 <= 4'h7; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_12 <= 4'h6;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_13 <= 4'h6; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_13 <= 4'h7;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_14 <= 4'hf; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_14 <= 4'he;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_15 <= 4'he; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_15 <= 4'hf;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_reg_data_r = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  out_reg_data_r_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  out_reg_data_r_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  out_reg_data_r_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  out_reg_data_r_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  out_reg_data_r_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  out_reg_data_r_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  out_reg_data_r_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  out_reg_data_r_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  out_reg_data_r_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  out_reg_data_r_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  out_reg_data_r_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  out_reg_data_r_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  out_reg_data_r_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  out_reg_data_r_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  out_reg_data_r_15 = _RAND_15[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Permute_switch_w16_bw64(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_0,
  input  [63:0] io_in_1,
  input  [63:0] io_in_2,
  input  [63:0] io_in_3,
  input  [63:0] io_in_4,
  input  [63:0] io_in_5,
  input  [63:0] io_in_6,
  input  [63:0] io_in_7,
  input  [63:0] io_in_8,
  input  [63:0] io_in_9,
  input  [63:0] io_in_10,
  input  [63:0] io_in_11,
  input  [63:0] io_in_12,
  input  [63:0] io_in_13,
  input  [63:0] io_in_14,
  input  [63:0] io_in_15,
  input  [3:0]  io_in_config_0,
  input  [3:0]  io_in_config_1,
  input  [3:0]  io_in_config_2,
  input  [3:0]  io_in_config_3,
  input  [3:0]  io_in_config_4,
  input  [3:0]  io_in_config_5,
  input  [3:0]  io_in_config_6,
  input  [3:0]  io_in_config_7,
  input  [3:0]  io_in_config_8,
  input  [3:0]  io_in_config_9,
  input  [3:0]  io_in_config_10,
  input  [3:0]  io_in_config_11,
  input  [3:0]  io_in_config_12,
  input  [3:0]  io_in_config_13,
  input  [3:0]  io_in_config_14,
  input  [3:0]  io_in_config_15,
  input         io_in_en,
  output        io_out_valid,
  output [63:0] io_out_0,
  output [63:0] io_out_1,
  output [63:0] io_out_2,
  output [63:0] io_out_3,
  output [63:0] io_out_4,
  output [63:0] io_out_5,
  output [63:0] io_out_6,
  output [63:0] io_out_7,
  output [63:0] io_out_8,
  output [63:0] io_out_9,
  output [63:0] io_out_10,
  output [63:0] io_out_11,
  output [63:0] io_out_12,
  output [63:0] io_out_13,
  output [63:0] io_out_14,
  output [63:0] io_out_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] dout_0; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_1; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_2; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_3; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_4; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_5; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_6; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_7; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_8; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_9; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_10; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_11; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_12; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_13; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_14; // @[PermutationDesigns.scala 198:23]
  reg [63:0] dout_15; // @[PermutationDesigns.scala 198:23]
  wire [63:0] _GEN_0 = 4'h0 == io_in_config_0 ? io_in_0 : dout_0; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_1 = 4'h1 == io_in_config_0 ? io_in_0 : dout_1; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_2 = 4'h2 == io_in_config_0 ? io_in_0 : dout_2; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_3 = 4'h3 == io_in_config_0 ? io_in_0 : dout_3; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_4 = 4'h4 == io_in_config_0 ? io_in_0 : dout_4; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_5 = 4'h5 == io_in_config_0 ? io_in_0 : dout_5; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_6 = 4'h6 == io_in_config_0 ? io_in_0 : dout_6; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_7 = 4'h7 == io_in_config_0 ? io_in_0 : dout_7; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_8 = 4'h8 == io_in_config_0 ? io_in_0 : dout_8; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_9 = 4'h9 == io_in_config_0 ? io_in_0 : dout_9; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_10 = 4'ha == io_in_config_0 ? io_in_0 : dout_10; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_11 = 4'hb == io_in_config_0 ? io_in_0 : dout_11; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_12 = 4'hc == io_in_config_0 ? io_in_0 : dout_12; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_13 = 4'hd == io_in_config_0 ? io_in_0 : dout_13; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_14 = 4'he == io_in_config_0 ? io_in_0 : dout_14; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_15 = 4'hf == io_in_config_0 ? io_in_0 : dout_15; // @[PermutationDesigns.scala 198:23 201:{31,31}]
  wire [63:0] _GEN_16 = io_in_en ? _GEN_0 : dout_0; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_17 = io_in_en ? _GEN_1 : dout_1; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_18 = io_in_en ? _GEN_2 : dout_2; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_19 = io_in_en ? _GEN_3 : dout_3; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_20 = io_in_en ? _GEN_4 : dout_4; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_21 = io_in_en ? _GEN_5 : dout_5; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_22 = io_in_en ? _GEN_6 : dout_6; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_23 = io_in_en ? _GEN_7 : dout_7; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_24 = io_in_en ? _GEN_8 : dout_8; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_25 = io_in_en ? _GEN_9 : dout_9; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_26 = io_in_en ? _GEN_10 : dout_10; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_27 = io_in_en ? _GEN_11 : dout_11; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_28 = io_in_en ? _GEN_12 : dout_12; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_29 = io_in_en ? _GEN_13 : dout_13; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_30 = io_in_en ? _GEN_14 : dout_14; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_31 = io_in_en ? _GEN_15 : dout_15; // @[PermutationDesigns.scala 200:21 198:23]
  wire [63:0] _GEN_32 = 4'h0 == io_in_config_1 ? io_in_1 : _GEN_16; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_33 = 4'h1 == io_in_config_1 ? io_in_1 : _GEN_17; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_34 = 4'h2 == io_in_config_1 ? io_in_1 : _GEN_18; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_35 = 4'h3 == io_in_config_1 ? io_in_1 : _GEN_19; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_36 = 4'h4 == io_in_config_1 ? io_in_1 : _GEN_20; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_37 = 4'h5 == io_in_config_1 ? io_in_1 : _GEN_21; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_38 = 4'h6 == io_in_config_1 ? io_in_1 : _GEN_22; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_39 = 4'h7 == io_in_config_1 ? io_in_1 : _GEN_23; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_40 = 4'h8 == io_in_config_1 ? io_in_1 : _GEN_24; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_41 = 4'h9 == io_in_config_1 ? io_in_1 : _GEN_25; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_42 = 4'ha == io_in_config_1 ? io_in_1 : _GEN_26; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_43 = 4'hb == io_in_config_1 ? io_in_1 : _GEN_27; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_44 = 4'hc == io_in_config_1 ? io_in_1 : _GEN_28; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_45 = 4'hd == io_in_config_1 ? io_in_1 : _GEN_29; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_46 = 4'he == io_in_config_1 ? io_in_1 : _GEN_30; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_47 = 4'hf == io_in_config_1 ? io_in_1 : _GEN_31; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_48 = io_in_en ? _GEN_32 : _GEN_16; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_49 = io_in_en ? _GEN_33 : _GEN_17; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_50 = io_in_en ? _GEN_34 : _GEN_18; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_51 = io_in_en ? _GEN_35 : _GEN_19; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_52 = io_in_en ? _GEN_36 : _GEN_20; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_53 = io_in_en ? _GEN_37 : _GEN_21; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_54 = io_in_en ? _GEN_38 : _GEN_22; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_55 = io_in_en ? _GEN_39 : _GEN_23; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_56 = io_in_en ? _GEN_40 : _GEN_24; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_57 = io_in_en ? _GEN_41 : _GEN_25; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_58 = io_in_en ? _GEN_42 : _GEN_26; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_59 = io_in_en ? _GEN_43 : _GEN_27; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_60 = io_in_en ? _GEN_44 : _GEN_28; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_61 = io_in_en ? _GEN_45 : _GEN_29; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_62 = io_in_en ? _GEN_46 : _GEN_30; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_63 = io_in_en ? _GEN_47 : _GEN_31; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_64 = 4'h0 == io_in_config_2 ? io_in_2 : _GEN_48; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_65 = 4'h1 == io_in_config_2 ? io_in_2 : _GEN_49; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_66 = 4'h2 == io_in_config_2 ? io_in_2 : _GEN_50; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_67 = 4'h3 == io_in_config_2 ? io_in_2 : _GEN_51; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_68 = 4'h4 == io_in_config_2 ? io_in_2 : _GEN_52; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_69 = 4'h5 == io_in_config_2 ? io_in_2 : _GEN_53; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_70 = 4'h6 == io_in_config_2 ? io_in_2 : _GEN_54; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_71 = 4'h7 == io_in_config_2 ? io_in_2 : _GEN_55; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_72 = 4'h8 == io_in_config_2 ? io_in_2 : _GEN_56; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_73 = 4'h9 == io_in_config_2 ? io_in_2 : _GEN_57; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_74 = 4'ha == io_in_config_2 ? io_in_2 : _GEN_58; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_75 = 4'hb == io_in_config_2 ? io_in_2 : _GEN_59; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_76 = 4'hc == io_in_config_2 ? io_in_2 : _GEN_60; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_77 = 4'hd == io_in_config_2 ? io_in_2 : _GEN_61; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_78 = 4'he == io_in_config_2 ? io_in_2 : _GEN_62; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_79 = 4'hf == io_in_config_2 ? io_in_2 : _GEN_63; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_80 = io_in_en ? _GEN_64 : _GEN_48; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_81 = io_in_en ? _GEN_65 : _GEN_49; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_82 = io_in_en ? _GEN_66 : _GEN_50; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_83 = io_in_en ? _GEN_67 : _GEN_51; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_84 = io_in_en ? _GEN_68 : _GEN_52; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_85 = io_in_en ? _GEN_69 : _GEN_53; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_86 = io_in_en ? _GEN_70 : _GEN_54; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_87 = io_in_en ? _GEN_71 : _GEN_55; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_88 = io_in_en ? _GEN_72 : _GEN_56; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_89 = io_in_en ? _GEN_73 : _GEN_57; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_90 = io_in_en ? _GEN_74 : _GEN_58; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_91 = io_in_en ? _GEN_75 : _GEN_59; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_92 = io_in_en ? _GEN_76 : _GEN_60; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_93 = io_in_en ? _GEN_77 : _GEN_61; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_94 = io_in_en ? _GEN_78 : _GEN_62; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_95 = io_in_en ? _GEN_79 : _GEN_63; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_96 = 4'h0 == io_in_config_3 ? io_in_3 : _GEN_80; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_97 = 4'h1 == io_in_config_3 ? io_in_3 : _GEN_81; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_98 = 4'h2 == io_in_config_3 ? io_in_3 : _GEN_82; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_99 = 4'h3 == io_in_config_3 ? io_in_3 : _GEN_83; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_100 = 4'h4 == io_in_config_3 ? io_in_3 : _GEN_84; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_101 = 4'h5 == io_in_config_3 ? io_in_3 : _GEN_85; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_102 = 4'h6 == io_in_config_3 ? io_in_3 : _GEN_86; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_103 = 4'h7 == io_in_config_3 ? io_in_3 : _GEN_87; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_104 = 4'h8 == io_in_config_3 ? io_in_3 : _GEN_88; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_105 = 4'h9 == io_in_config_3 ? io_in_3 : _GEN_89; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_106 = 4'ha == io_in_config_3 ? io_in_3 : _GEN_90; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_107 = 4'hb == io_in_config_3 ? io_in_3 : _GEN_91; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_108 = 4'hc == io_in_config_3 ? io_in_3 : _GEN_92; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_109 = 4'hd == io_in_config_3 ? io_in_3 : _GEN_93; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_110 = 4'he == io_in_config_3 ? io_in_3 : _GEN_94; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_111 = 4'hf == io_in_config_3 ? io_in_3 : _GEN_95; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_112 = io_in_en ? _GEN_96 : _GEN_80; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_113 = io_in_en ? _GEN_97 : _GEN_81; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_114 = io_in_en ? _GEN_98 : _GEN_82; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_115 = io_in_en ? _GEN_99 : _GEN_83; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_116 = io_in_en ? _GEN_100 : _GEN_84; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_117 = io_in_en ? _GEN_101 : _GEN_85; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_118 = io_in_en ? _GEN_102 : _GEN_86; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_119 = io_in_en ? _GEN_103 : _GEN_87; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_120 = io_in_en ? _GEN_104 : _GEN_88; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_121 = io_in_en ? _GEN_105 : _GEN_89; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_122 = io_in_en ? _GEN_106 : _GEN_90; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_123 = io_in_en ? _GEN_107 : _GEN_91; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_124 = io_in_en ? _GEN_108 : _GEN_92; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_125 = io_in_en ? _GEN_109 : _GEN_93; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_126 = io_in_en ? _GEN_110 : _GEN_94; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_127 = io_in_en ? _GEN_111 : _GEN_95; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_128 = 4'h0 == io_in_config_4 ? io_in_4 : _GEN_112; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_129 = 4'h1 == io_in_config_4 ? io_in_4 : _GEN_113; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_130 = 4'h2 == io_in_config_4 ? io_in_4 : _GEN_114; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_131 = 4'h3 == io_in_config_4 ? io_in_4 : _GEN_115; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_132 = 4'h4 == io_in_config_4 ? io_in_4 : _GEN_116; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_133 = 4'h5 == io_in_config_4 ? io_in_4 : _GEN_117; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_134 = 4'h6 == io_in_config_4 ? io_in_4 : _GEN_118; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_135 = 4'h7 == io_in_config_4 ? io_in_4 : _GEN_119; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_136 = 4'h8 == io_in_config_4 ? io_in_4 : _GEN_120; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_137 = 4'h9 == io_in_config_4 ? io_in_4 : _GEN_121; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_138 = 4'ha == io_in_config_4 ? io_in_4 : _GEN_122; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_139 = 4'hb == io_in_config_4 ? io_in_4 : _GEN_123; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_140 = 4'hc == io_in_config_4 ? io_in_4 : _GEN_124; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_141 = 4'hd == io_in_config_4 ? io_in_4 : _GEN_125; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_142 = 4'he == io_in_config_4 ? io_in_4 : _GEN_126; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_143 = 4'hf == io_in_config_4 ? io_in_4 : _GEN_127; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_144 = io_in_en ? _GEN_128 : _GEN_112; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_145 = io_in_en ? _GEN_129 : _GEN_113; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_146 = io_in_en ? _GEN_130 : _GEN_114; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_147 = io_in_en ? _GEN_131 : _GEN_115; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_148 = io_in_en ? _GEN_132 : _GEN_116; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_149 = io_in_en ? _GEN_133 : _GEN_117; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_150 = io_in_en ? _GEN_134 : _GEN_118; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_151 = io_in_en ? _GEN_135 : _GEN_119; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_152 = io_in_en ? _GEN_136 : _GEN_120; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_153 = io_in_en ? _GEN_137 : _GEN_121; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_154 = io_in_en ? _GEN_138 : _GEN_122; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_155 = io_in_en ? _GEN_139 : _GEN_123; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_156 = io_in_en ? _GEN_140 : _GEN_124; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_157 = io_in_en ? _GEN_141 : _GEN_125; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_158 = io_in_en ? _GEN_142 : _GEN_126; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_159 = io_in_en ? _GEN_143 : _GEN_127; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_160 = 4'h0 == io_in_config_5 ? io_in_5 : _GEN_144; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_161 = 4'h1 == io_in_config_5 ? io_in_5 : _GEN_145; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_162 = 4'h2 == io_in_config_5 ? io_in_5 : _GEN_146; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_163 = 4'h3 == io_in_config_5 ? io_in_5 : _GEN_147; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_164 = 4'h4 == io_in_config_5 ? io_in_5 : _GEN_148; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_165 = 4'h5 == io_in_config_5 ? io_in_5 : _GEN_149; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_166 = 4'h6 == io_in_config_5 ? io_in_5 : _GEN_150; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_167 = 4'h7 == io_in_config_5 ? io_in_5 : _GEN_151; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_168 = 4'h8 == io_in_config_5 ? io_in_5 : _GEN_152; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_169 = 4'h9 == io_in_config_5 ? io_in_5 : _GEN_153; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_170 = 4'ha == io_in_config_5 ? io_in_5 : _GEN_154; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_171 = 4'hb == io_in_config_5 ? io_in_5 : _GEN_155; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_172 = 4'hc == io_in_config_5 ? io_in_5 : _GEN_156; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_173 = 4'hd == io_in_config_5 ? io_in_5 : _GEN_157; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_174 = 4'he == io_in_config_5 ? io_in_5 : _GEN_158; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_175 = 4'hf == io_in_config_5 ? io_in_5 : _GEN_159; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_176 = io_in_en ? _GEN_160 : _GEN_144; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_177 = io_in_en ? _GEN_161 : _GEN_145; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_178 = io_in_en ? _GEN_162 : _GEN_146; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_179 = io_in_en ? _GEN_163 : _GEN_147; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_180 = io_in_en ? _GEN_164 : _GEN_148; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_181 = io_in_en ? _GEN_165 : _GEN_149; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_182 = io_in_en ? _GEN_166 : _GEN_150; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_183 = io_in_en ? _GEN_167 : _GEN_151; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_184 = io_in_en ? _GEN_168 : _GEN_152; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_185 = io_in_en ? _GEN_169 : _GEN_153; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_186 = io_in_en ? _GEN_170 : _GEN_154; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_187 = io_in_en ? _GEN_171 : _GEN_155; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_188 = io_in_en ? _GEN_172 : _GEN_156; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_189 = io_in_en ? _GEN_173 : _GEN_157; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_190 = io_in_en ? _GEN_174 : _GEN_158; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_191 = io_in_en ? _GEN_175 : _GEN_159; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_192 = 4'h0 == io_in_config_6 ? io_in_6 : _GEN_176; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_193 = 4'h1 == io_in_config_6 ? io_in_6 : _GEN_177; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_194 = 4'h2 == io_in_config_6 ? io_in_6 : _GEN_178; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_195 = 4'h3 == io_in_config_6 ? io_in_6 : _GEN_179; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_196 = 4'h4 == io_in_config_6 ? io_in_6 : _GEN_180; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_197 = 4'h5 == io_in_config_6 ? io_in_6 : _GEN_181; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_198 = 4'h6 == io_in_config_6 ? io_in_6 : _GEN_182; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_199 = 4'h7 == io_in_config_6 ? io_in_6 : _GEN_183; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_200 = 4'h8 == io_in_config_6 ? io_in_6 : _GEN_184; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_201 = 4'h9 == io_in_config_6 ? io_in_6 : _GEN_185; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_202 = 4'ha == io_in_config_6 ? io_in_6 : _GEN_186; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_203 = 4'hb == io_in_config_6 ? io_in_6 : _GEN_187; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_204 = 4'hc == io_in_config_6 ? io_in_6 : _GEN_188; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_205 = 4'hd == io_in_config_6 ? io_in_6 : _GEN_189; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_206 = 4'he == io_in_config_6 ? io_in_6 : _GEN_190; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_207 = 4'hf == io_in_config_6 ? io_in_6 : _GEN_191; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_208 = io_in_en ? _GEN_192 : _GEN_176; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_209 = io_in_en ? _GEN_193 : _GEN_177; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_210 = io_in_en ? _GEN_194 : _GEN_178; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_211 = io_in_en ? _GEN_195 : _GEN_179; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_212 = io_in_en ? _GEN_196 : _GEN_180; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_213 = io_in_en ? _GEN_197 : _GEN_181; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_214 = io_in_en ? _GEN_198 : _GEN_182; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_215 = io_in_en ? _GEN_199 : _GEN_183; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_216 = io_in_en ? _GEN_200 : _GEN_184; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_217 = io_in_en ? _GEN_201 : _GEN_185; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_218 = io_in_en ? _GEN_202 : _GEN_186; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_219 = io_in_en ? _GEN_203 : _GEN_187; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_220 = io_in_en ? _GEN_204 : _GEN_188; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_221 = io_in_en ? _GEN_205 : _GEN_189; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_222 = io_in_en ? _GEN_206 : _GEN_190; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_223 = io_in_en ? _GEN_207 : _GEN_191; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_224 = 4'h0 == io_in_config_7 ? io_in_7 : _GEN_208; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_225 = 4'h1 == io_in_config_7 ? io_in_7 : _GEN_209; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_226 = 4'h2 == io_in_config_7 ? io_in_7 : _GEN_210; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_227 = 4'h3 == io_in_config_7 ? io_in_7 : _GEN_211; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_228 = 4'h4 == io_in_config_7 ? io_in_7 : _GEN_212; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_229 = 4'h5 == io_in_config_7 ? io_in_7 : _GEN_213; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_230 = 4'h6 == io_in_config_7 ? io_in_7 : _GEN_214; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_231 = 4'h7 == io_in_config_7 ? io_in_7 : _GEN_215; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_232 = 4'h8 == io_in_config_7 ? io_in_7 : _GEN_216; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_233 = 4'h9 == io_in_config_7 ? io_in_7 : _GEN_217; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_234 = 4'ha == io_in_config_7 ? io_in_7 : _GEN_218; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_235 = 4'hb == io_in_config_7 ? io_in_7 : _GEN_219; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_236 = 4'hc == io_in_config_7 ? io_in_7 : _GEN_220; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_237 = 4'hd == io_in_config_7 ? io_in_7 : _GEN_221; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_238 = 4'he == io_in_config_7 ? io_in_7 : _GEN_222; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_239 = 4'hf == io_in_config_7 ? io_in_7 : _GEN_223; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_240 = io_in_en ? _GEN_224 : _GEN_208; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_241 = io_in_en ? _GEN_225 : _GEN_209; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_242 = io_in_en ? _GEN_226 : _GEN_210; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_243 = io_in_en ? _GEN_227 : _GEN_211; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_244 = io_in_en ? _GEN_228 : _GEN_212; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_245 = io_in_en ? _GEN_229 : _GEN_213; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_246 = io_in_en ? _GEN_230 : _GEN_214; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_247 = io_in_en ? _GEN_231 : _GEN_215; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_248 = io_in_en ? _GEN_232 : _GEN_216; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_249 = io_in_en ? _GEN_233 : _GEN_217; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_250 = io_in_en ? _GEN_234 : _GEN_218; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_251 = io_in_en ? _GEN_235 : _GEN_219; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_252 = io_in_en ? _GEN_236 : _GEN_220; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_253 = io_in_en ? _GEN_237 : _GEN_221; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_254 = io_in_en ? _GEN_238 : _GEN_222; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_255 = io_in_en ? _GEN_239 : _GEN_223; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_256 = 4'h0 == io_in_config_8 ? io_in_8 : _GEN_240; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_257 = 4'h1 == io_in_config_8 ? io_in_8 : _GEN_241; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_258 = 4'h2 == io_in_config_8 ? io_in_8 : _GEN_242; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_259 = 4'h3 == io_in_config_8 ? io_in_8 : _GEN_243; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_260 = 4'h4 == io_in_config_8 ? io_in_8 : _GEN_244; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_261 = 4'h5 == io_in_config_8 ? io_in_8 : _GEN_245; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_262 = 4'h6 == io_in_config_8 ? io_in_8 : _GEN_246; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_263 = 4'h7 == io_in_config_8 ? io_in_8 : _GEN_247; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_264 = 4'h8 == io_in_config_8 ? io_in_8 : _GEN_248; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_265 = 4'h9 == io_in_config_8 ? io_in_8 : _GEN_249; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_266 = 4'ha == io_in_config_8 ? io_in_8 : _GEN_250; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_267 = 4'hb == io_in_config_8 ? io_in_8 : _GEN_251; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_268 = 4'hc == io_in_config_8 ? io_in_8 : _GEN_252; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_269 = 4'hd == io_in_config_8 ? io_in_8 : _GEN_253; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_270 = 4'he == io_in_config_8 ? io_in_8 : _GEN_254; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_271 = 4'hf == io_in_config_8 ? io_in_8 : _GEN_255; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_272 = io_in_en ? _GEN_256 : _GEN_240; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_273 = io_in_en ? _GEN_257 : _GEN_241; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_274 = io_in_en ? _GEN_258 : _GEN_242; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_275 = io_in_en ? _GEN_259 : _GEN_243; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_276 = io_in_en ? _GEN_260 : _GEN_244; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_277 = io_in_en ? _GEN_261 : _GEN_245; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_278 = io_in_en ? _GEN_262 : _GEN_246; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_279 = io_in_en ? _GEN_263 : _GEN_247; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_280 = io_in_en ? _GEN_264 : _GEN_248; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_281 = io_in_en ? _GEN_265 : _GEN_249; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_282 = io_in_en ? _GEN_266 : _GEN_250; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_283 = io_in_en ? _GEN_267 : _GEN_251; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_284 = io_in_en ? _GEN_268 : _GEN_252; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_285 = io_in_en ? _GEN_269 : _GEN_253; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_286 = io_in_en ? _GEN_270 : _GEN_254; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_287 = io_in_en ? _GEN_271 : _GEN_255; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_288 = 4'h0 == io_in_config_9 ? io_in_9 : _GEN_272; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_289 = 4'h1 == io_in_config_9 ? io_in_9 : _GEN_273; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_290 = 4'h2 == io_in_config_9 ? io_in_9 : _GEN_274; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_291 = 4'h3 == io_in_config_9 ? io_in_9 : _GEN_275; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_292 = 4'h4 == io_in_config_9 ? io_in_9 : _GEN_276; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_293 = 4'h5 == io_in_config_9 ? io_in_9 : _GEN_277; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_294 = 4'h6 == io_in_config_9 ? io_in_9 : _GEN_278; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_295 = 4'h7 == io_in_config_9 ? io_in_9 : _GEN_279; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_296 = 4'h8 == io_in_config_9 ? io_in_9 : _GEN_280; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_297 = 4'h9 == io_in_config_9 ? io_in_9 : _GEN_281; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_298 = 4'ha == io_in_config_9 ? io_in_9 : _GEN_282; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_299 = 4'hb == io_in_config_9 ? io_in_9 : _GEN_283; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_300 = 4'hc == io_in_config_9 ? io_in_9 : _GEN_284; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_301 = 4'hd == io_in_config_9 ? io_in_9 : _GEN_285; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_302 = 4'he == io_in_config_9 ? io_in_9 : _GEN_286; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_303 = 4'hf == io_in_config_9 ? io_in_9 : _GEN_287; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_304 = io_in_en ? _GEN_288 : _GEN_272; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_305 = io_in_en ? _GEN_289 : _GEN_273; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_306 = io_in_en ? _GEN_290 : _GEN_274; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_307 = io_in_en ? _GEN_291 : _GEN_275; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_308 = io_in_en ? _GEN_292 : _GEN_276; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_309 = io_in_en ? _GEN_293 : _GEN_277; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_310 = io_in_en ? _GEN_294 : _GEN_278; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_311 = io_in_en ? _GEN_295 : _GEN_279; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_312 = io_in_en ? _GEN_296 : _GEN_280; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_313 = io_in_en ? _GEN_297 : _GEN_281; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_314 = io_in_en ? _GEN_298 : _GEN_282; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_315 = io_in_en ? _GEN_299 : _GEN_283; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_316 = io_in_en ? _GEN_300 : _GEN_284; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_317 = io_in_en ? _GEN_301 : _GEN_285; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_318 = io_in_en ? _GEN_302 : _GEN_286; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_319 = io_in_en ? _GEN_303 : _GEN_287; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_320 = 4'h0 == io_in_config_10 ? io_in_10 : _GEN_304; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_321 = 4'h1 == io_in_config_10 ? io_in_10 : _GEN_305; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_322 = 4'h2 == io_in_config_10 ? io_in_10 : _GEN_306; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_323 = 4'h3 == io_in_config_10 ? io_in_10 : _GEN_307; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_324 = 4'h4 == io_in_config_10 ? io_in_10 : _GEN_308; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_325 = 4'h5 == io_in_config_10 ? io_in_10 : _GEN_309; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_326 = 4'h6 == io_in_config_10 ? io_in_10 : _GEN_310; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_327 = 4'h7 == io_in_config_10 ? io_in_10 : _GEN_311; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_328 = 4'h8 == io_in_config_10 ? io_in_10 : _GEN_312; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_329 = 4'h9 == io_in_config_10 ? io_in_10 : _GEN_313; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_330 = 4'ha == io_in_config_10 ? io_in_10 : _GEN_314; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_331 = 4'hb == io_in_config_10 ? io_in_10 : _GEN_315; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_332 = 4'hc == io_in_config_10 ? io_in_10 : _GEN_316; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_333 = 4'hd == io_in_config_10 ? io_in_10 : _GEN_317; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_334 = 4'he == io_in_config_10 ? io_in_10 : _GEN_318; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_335 = 4'hf == io_in_config_10 ? io_in_10 : _GEN_319; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_336 = io_in_en ? _GEN_320 : _GEN_304; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_337 = io_in_en ? _GEN_321 : _GEN_305; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_338 = io_in_en ? _GEN_322 : _GEN_306; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_339 = io_in_en ? _GEN_323 : _GEN_307; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_340 = io_in_en ? _GEN_324 : _GEN_308; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_341 = io_in_en ? _GEN_325 : _GEN_309; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_342 = io_in_en ? _GEN_326 : _GEN_310; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_343 = io_in_en ? _GEN_327 : _GEN_311; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_344 = io_in_en ? _GEN_328 : _GEN_312; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_345 = io_in_en ? _GEN_329 : _GEN_313; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_346 = io_in_en ? _GEN_330 : _GEN_314; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_347 = io_in_en ? _GEN_331 : _GEN_315; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_348 = io_in_en ? _GEN_332 : _GEN_316; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_349 = io_in_en ? _GEN_333 : _GEN_317; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_350 = io_in_en ? _GEN_334 : _GEN_318; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_351 = io_in_en ? _GEN_335 : _GEN_319; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_352 = 4'h0 == io_in_config_11 ? io_in_11 : _GEN_336; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_353 = 4'h1 == io_in_config_11 ? io_in_11 : _GEN_337; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_354 = 4'h2 == io_in_config_11 ? io_in_11 : _GEN_338; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_355 = 4'h3 == io_in_config_11 ? io_in_11 : _GEN_339; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_356 = 4'h4 == io_in_config_11 ? io_in_11 : _GEN_340; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_357 = 4'h5 == io_in_config_11 ? io_in_11 : _GEN_341; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_358 = 4'h6 == io_in_config_11 ? io_in_11 : _GEN_342; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_359 = 4'h7 == io_in_config_11 ? io_in_11 : _GEN_343; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_360 = 4'h8 == io_in_config_11 ? io_in_11 : _GEN_344; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_361 = 4'h9 == io_in_config_11 ? io_in_11 : _GEN_345; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_362 = 4'ha == io_in_config_11 ? io_in_11 : _GEN_346; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_363 = 4'hb == io_in_config_11 ? io_in_11 : _GEN_347; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_364 = 4'hc == io_in_config_11 ? io_in_11 : _GEN_348; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_365 = 4'hd == io_in_config_11 ? io_in_11 : _GEN_349; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_366 = 4'he == io_in_config_11 ? io_in_11 : _GEN_350; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_367 = 4'hf == io_in_config_11 ? io_in_11 : _GEN_351; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_368 = io_in_en ? _GEN_352 : _GEN_336; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_369 = io_in_en ? _GEN_353 : _GEN_337; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_370 = io_in_en ? _GEN_354 : _GEN_338; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_371 = io_in_en ? _GEN_355 : _GEN_339; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_372 = io_in_en ? _GEN_356 : _GEN_340; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_373 = io_in_en ? _GEN_357 : _GEN_341; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_374 = io_in_en ? _GEN_358 : _GEN_342; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_375 = io_in_en ? _GEN_359 : _GEN_343; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_376 = io_in_en ? _GEN_360 : _GEN_344; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_377 = io_in_en ? _GEN_361 : _GEN_345; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_378 = io_in_en ? _GEN_362 : _GEN_346; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_379 = io_in_en ? _GEN_363 : _GEN_347; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_380 = io_in_en ? _GEN_364 : _GEN_348; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_381 = io_in_en ? _GEN_365 : _GEN_349; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_382 = io_in_en ? _GEN_366 : _GEN_350; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_383 = io_in_en ? _GEN_367 : _GEN_351; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_384 = 4'h0 == io_in_config_12 ? io_in_12 : _GEN_368; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_385 = 4'h1 == io_in_config_12 ? io_in_12 : _GEN_369; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_386 = 4'h2 == io_in_config_12 ? io_in_12 : _GEN_370; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_387 = 4'h3 == io_in_config_12 ? io_in_12 : _GEN_371; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_388 = 4'h4 == io_in_config_12 ? io_in_12 : _GEN_372; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_389 = 4'h5 == io_in_config_12 ? io_in_12 : _GEN_373; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_390 = 4'h6 == io_in_config_12 ? io_in_12 : _GEN_374; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_391 = 4'h7 == io_in_config_12 ? io_in_12 : _GEN_375; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_392 = 4'h8 == io_in_config_12 ? io_in_12 : _GEN_376; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_393 = 4'h9 == io_in_config_12 ? io_in_12 : _GEN_377; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_394 = 4'ha == io_in_config_12 ? io_in_12 : _GEN_378; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_395 = 4'hb == io_in_config_12 ? io_in_12 : _GEN_379; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_396 = 4'hc == io_in_config_12 ? io_in_12 : _GEN_380; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_397 = 4'hd == io_in_config_12 ? io_in_12 : _GEN_381; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_398 = 4'he == io_in_config_12 ? io_in_12 : _GEN_382; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_399 = 4'hf == io_in_config_12 ? io_in_12 : _GEN_383; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_400 = io_in_en ? _GEN_384 : _GEN_368; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_401 = io_in_en ? _GEN_385 : _GEN_369; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_402 = io_in_en ? _GEN_386 : _GEN_370; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_403 = io_in_en ? _GEN_387 : _GEN_371; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_404 = io_in_en ? _GEN_388 : _GEN_372; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_405 = io_in_en ? _GEN_389 : _GEN_373; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_406 = io_in_en ? _GEN_390 : _GEN_374; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_407 = io_in_en ? _GEN_391 : _GEN_375; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_408 = io_in_en ? _GEN_392 : _GEN_376; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_409 = io_in_en ? _GEN_393 : _GEN_377; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_410 = io_in_en ? _GEN_394 : _GEN_378; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_411 = io_in_en ? _GEN_395 : _GEN_379; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_412 = io_in_en ? _GEN_396 : _GEN_380; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_413 = io_in_en ? _GEN_397 : _GEN_381; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_414 = io_in_en ? _GEN_398 : _GEN_382; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_415 = io_in_en ? _GEN_399 : _GEN_383; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_416 = 4'h0 == io_in_config_13 ? io_in_13 : _GEN_400; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_417 = 4'h1 == io_in_config_13 ? io_in_13 : _GEN_401; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_418 = 4'h2 == io_in_config_13 ? io_in_13 : _GEN_402; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_419 = 4'h3 == io_in_config_13 ? io_in_13 : _GEN_403; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_420 = 4'h4 == io_in_config_13 ? io_in_13 : _GEN_404; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_421 = 4'h5 == io_in_config_13 ? io_in_13 : _GEN_405; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_422 = 4'h6 == io_in_config_13 ? io_in_13 : _GEN_406; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_423 = 4'h7 == io_in_config_13 ? io_in_13 : _GEN_407; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_424 = 4'h8 == io_in_config_13 ? io_in_13 : _GEN_408; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_425 = 4'h9 == io_in_config_13 ? io_in_13 : _GEN_409; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_426 = 4'ha == io_in_config_13 ? io_in_13 : _GEN_410; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_427 = 4'hb == io_in_config_13 ? io_in_13 : _GEN_411; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_428 = 4'hc == io_in_config_13 ? io_in_13 : _GEN_412; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_429 = 4'hd == io_in_config_13 ? io_in_13 : _GEN_413; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_430 = 4'he == io_in_config_13 ? io_in_13 : _GEN_414; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_431 = 4'hf == io_in_config_13 ? io_in_13 : _GEN_415; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_432 = io_in_en ? _GEN_416 : _GEN_400; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_433 = io_in_en ? _GEN_417 : _GEN_401; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_434 = io_in_en ? _GEN_418 : _GEN_402; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_435 = io_in_en ? _GEN_419 : _GEN_403; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_436 = io_in_en ? _GEN_420 : _GEN_404; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_437 = io_in_en ? _GEN_421 : _GEN_405; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_438 = io_in_en ? _GEN_422 : _GEN_406; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_439 = io_in_en ? _GEN_423 : _GEN_407; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_440 = io_in_en ? _GEN_424 : _GEN_408; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_441 = io_in_en ? _GEN_425 : _GEN_409; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_442 = io_in_en ? _GEN_426 : _GEN_410; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_443 = io_in_en ? _GEN_427 : _GEN_411; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_444 = io_in_en ? _GEN_428 : _GEN_412; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_445 = io_in_en ? _GEN_429 : _GEN_413; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_446 = io_in_en ? _GEN_430 : _GEN_414; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_447 = io_in_en ? _GEN_431 : _GEN_415; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_448 = 4'h0 == io_in_config_14 ? io_in_14 : _GEN_432; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_449 = 4'h1 == io_in_config_14 ? io_in_14 : _GEN_433; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_450 = 4'h2 == io_in_config_14 ? io_in_14 : _GEN_434; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_451 = 4'h3 == io_in_config_14 ? io_in_14 : _GEN_435; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_452 = 4'h4 == io_in_config_14 ? io_in_14 : _GEN_436; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_453 = 4'h5 == io_in_config_14 ? io_in_14 : _GEN_437; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_454 = 4'h6 == io_in_config_14 ? io_in_14 : _GEN_438; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_455 = 4'h7 == io_in_config_14 ? io_in_14 : _GEN_439; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_456 = 4'h8 == io_in_config_14 ? io_in_14 : _GEN_440; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_457 = 4'h9 == io_in_config_14 ? io_in_14 : _GEN_441; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_458 = 4'ha == io_in_config_14 ? io_in_14 : _GEN_442; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_459 = 4'hb == io_in_config_14 ? io_in_14 : _GEN_443; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_460 = 4'hc == io_in_config_14 ? io_in_14 : _GEN_444; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_461 = 4'hd == io_in_config_14 ? io_in_14 : _GEN_445; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_462 = 4'he == io_in_config_14 ? io_in_14 : _GEN_446; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_463 = 4'hf == io_in_config_14 ? io_in_14 : _GEN_447; // @[PermutationDesigns.scala 201:{31,31}]
  wire [63:0] _GEN_464 = io_in_en ? _GEN_448 : _GEN_432; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_465 = io_in_en ? _GEN_449 : _GEN_433; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_466 = io_in_en ? _GEN_450 : _GEN_434; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_467 = io_in_en ? _GEN_451 : _GEN_435; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_468 = io_in_en ? _GEN_452 : _GEN_436; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_469 = io_in_en ? _GEN_453 : _GEN_437; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_470 = io_in_en ? _GEN_454 : _GEN_438; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_471 = io_in_en ? _GEN_455 : _GEN_439; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_472 = io_in_en ? _GEN_456 : _GEN_440; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_473 = io_in_en ? _GEN_457 : _GEN_441; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_474 = io_in_en ? _GEN_458 : _GEN_442; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_475 = io_in_en ? _GEN_459 : _GEN_443; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_476 = io_in_en ? _GEN_460 : _GEN_444; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_477 = io_in_en ? _GEN_461 : _GEN_445; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_478 = io_in_en ? _GEN_462 : _GEN_446; // @[PermutationDesigns.scala 200:21]
  wire [63:0] _GEN_479 = io_in_en ? _GEN_463 : _GEN_447; // @[PermutationDesigns.scala 200:21]
  reg  io_out_valid_r; // @[Reg.scala 16:16]
  assign io_out_valid = io_out_valid_r; // @[PermutationDesigns.scala 205:18]
  assign io_out_0 = dout_0; // @[PermutationDesigns.scala 204:12]
  assign io_out_1 = dout_1; // @[PermutationDesigns.scala 204:12]
  assign io_out_2 = dout_2; // @[PermutationDesigns.scala 204:12]
  assign io_out_3 = dout_3; // @[PermutationDesigns.scala 204:12]
  assign io_out_4 = dout_4; // @[PermutationDesigns.scala 204:12]
  assign io_out_5 = dout_5; // @[PermutationDesigns.scala 204:12]
  assign io_out_6 = dout_6; // @[PermutationDesigns.scala 204:12]
  assign io_out_7 = dout_7; // @[PermutationDesigns.scala 204:12]
  assign io_out_8 = dout_8; // @[PermutationDesigns.scala 204:12]
  assign io_out_9 = dout_9; // @[PermutationDesigns.scala 204:12]
  assign io_out_10 = dout_10; // @[PermutationDesigns.scala 204:12]
  assign io_out_11 = dout_11; // @[PermutationDesigns.scala 204:12]
  assign io_out_12 = dout_12; // @[PermutationDesigns.scala 204:12]
  assign io_out_13 = dout_13; // @[PermutationDesigns.scala 204:12]
  assign io_out_14 = dout_14; // @[PermutationDesigns.scala 204:12]
  assign io_out_15 = dout_15; // @[PermutationDesigns.scala 204:12]
  always @(posedge clock) begin
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_0 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'h0 == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_0 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_0 <= _GEN_464;
      end
    end else begin
      dout_0 <= _GEN_464;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_1 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'h1 == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_1 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_1 <= _GEN_465;
      end
    end else begin
      dout_1 <= _GEN_465;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_2 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'h2 == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_2 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_2 <= _GEN_466;
      end
    end else begin
      dout_2 <= _GEN_466;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_3 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'h3 == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_3 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_3 <= _GEN_467;
      end
    end else begin
      dout_3 <= _GEN_467;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_4 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'h4 == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_4 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_4 <= _GEN_468;
      end
    end else begin
      dout_4 <= _GEN_468;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_5 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'h5 == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_5 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_5 <= _GEN_469;
      end
    end else begin
      dout_5 <= _GEN_469;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_6 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'h6 == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_6 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_6 <= _GEN_470;
      end
    end else begin
      dout_6 <= _GEN_470;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_7 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'h7 == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_7 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_7 <= _GEN_471;
      end
    end else begin
      dout_7 <= _GEN_471;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_8 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'h8 == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_8 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_8 <= _GEN_472;
      end
    end else begin
      dout_8 <= _GEN_472;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_9 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'h9 == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_9 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_9 <= _GEN_473;
      end
    end else begin
      dout_9 <= _GEN_473;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_10 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'ha == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_10 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_10 <= _GEN_474;
      end
    end else begin
      dout_10 <= _GEN_474;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_11 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'hb == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_11 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_11 <= _GEN_475;
      end
    end else begin
      dout_11 <= _GEN_475;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_12 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'hc == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_12 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_12 <= _GEN_476;
      end
    end else begin
      dout_12 <= _GEN_476;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_13 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'hd == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_13 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_13 <= _GEN_477;
      end
    end else begin
      dout_13 <= _GEN_477;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_14 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'he == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_14 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_14 <= _GEN_478;
      end
    end else begin
      dout_14 <= _GEN_478;
    end
    if (reset) begin // @[PermutationDesigns.scala 198:23]
      dout_15 <= 64'h0; // @[PermutationDesigns.scala 198:23]
    end else if (io_in_en) begin // @[PermutationDesigns.scala 200:21]
      if (4'hf == io_in_config_15) begin // @[PermutationDesigns.scala 201:31]
        dout_15 <= io_in_15; // @[PermutationDesigns.scala 201:31]
      end else begin
        dout_15 <= _GEN_479;
      end
    end else begin
      dout_15 <= _GEN_479;
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r <= io_in_valid; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  dout_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  dout_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  dout_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  dout_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  dout_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  dout_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dout_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dout_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dout_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  dout_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  dout_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  dout_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  dout_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  dout_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  dout_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  dout_15 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  io_out_valid_r = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2(
  input   clock,
  input   io_in_en,
  input   io_in_cnt,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg  out_reg_data_r; // @[Reg.scala 16:16]
  reg  out_reg_data_r_1; // @[Reg.scala 16:16]
  reg  out_reg_data_r_2; // @[Reg.scala 16:16]
  reg  out_reg_data_r_3; // @[Reg.scala 16:16]
  reg  out_reg_data_r_4; // @[Reg.scala 16:16]
  reg  out_reg_data_r_5; // @[Reg.scala 16:16]
  reg  out_reg_data_r_6; // @[Reg.scala 16:16]
  reg  out_reg_data_r_7; // @[Reg.scala 16:16]
  reg  out_reg_data_r_8; // @[Reg.scala 16:16]
  reg  out_reg_data_r_9; // @[Reg.scala 16:16]
  reg  out_reg_data_r_10; // @[Reg.scala 16:16]
  reg  out_reg_data_r_11; // @[Reg.scala 16:16]
  reg  out_reg_data_r_12; // @[Reg.scala 16:16]
  reg  out_reg_data_r_13; // @[Reg.scala 16:16]
  reg  out_reg_data_r_14; // @[Reg.scala 16:16]
  reg  out_reg_data_r_15; // @[Reg.scala 16:16]
  assign io_out_0 = out_reg_data_r; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_1 = out_reg_data_r_1; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_2 = out_reg_data_r_2; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_3 = out_reg_data_r_3; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_4 = out_reg_data_r_4; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_5 = out_reg_data_r_5; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_6 = out_reg_data_r_6; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_7 = out_reg_data_r_7; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_8 = out_reg_data_r_8; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_9 = out_reg_data_r_9; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_10 = out_reg_data_r_10; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_11 = out_reg_data_r_11; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_12 = out_reg_data_r_12; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_13 = out_reg_data_r_13; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_14 = out_reg_data_r_14; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_15 = out_reg_data_r_15; // @[PermutationDesigns.scala 229:{31,31}]
  always @(posedge clock) begin
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_1 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_1 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_2 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_3 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_3 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_4 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_5 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_5 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_6 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_7 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_7 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_8 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_9 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_9 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_10 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_11 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_11 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_12 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_13 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_13 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_14 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_15 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_15 <= 1'h1;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_reg_data_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_reg_data_r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_reg_data_r_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_reg_data_r_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_reg_data_r_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_reg_data_r_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_reg_data_r_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  out_reg_data_r_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  out_reg_data_r_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  out_reg_data_r_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  out_reg_data_r_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  out_reg_data_r_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  out_reg_data_r_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  out_reg_data_r_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  out_reg_data_r_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  out_reg_data_r_15 = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Permute_Streaming_N32_r2_w16_bitRtrue_bw64(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [63:0] io_in_0,
  input  [63:0] io_in_1,
  input  [63:0] io_in_2,
  input  [63:0] io_in_3,
  input  [63:0] io_in_4,
  input  [63:0] io_in_5,
  input  [63:0] io_in_6,
  input  [63:0] io_in_7,
  input  [63:0] io_in_8,
  input  [63:0] io_in_9,
  input  [63:0] io_in_10,
  input  [63:0] io_in_11,
  input  [63:0] io_in_12,
  input  [63:0] io_in_13,
  input  [63:0] io_in_14,
  input  [63:0] io_in_15,
  input         io_in_valid,
  output [63:0] io_out_0,
  output [63:0] io_out_1,
  output [63:0] io_out_2,
  output [63:0] io_out_3,
  output [63:0] io_out_4,
  output [63:0] io_out_5,
  output [63:0] io_out_6,
  output [63:0] io_out_7,
  output [63:0] io_out_8,
  output [63:0] io_out_9,
  output [63:0] io_out_10,
  output [63:0] io_out_11,
  output [63:0] io_out_12,
  output [63:0] io_out_13,
  output [63:0] io_out_14,
  output [63:0] io_out_15,
  output        io_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_Block_N32_w16_bw64_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_1_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_1_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_1_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_1_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_1_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_1_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_1_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_1_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_2_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_2_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_2_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_2_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_2_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_2_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_2_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_2_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_3_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_3_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_3_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_3_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_3_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_3_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_3_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_3_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_4_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_4_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_4_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_4_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_4_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_4_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_4_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_4_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_5_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_5_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_5_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_5_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_5_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_5_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_5_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_5_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_6_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_6_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_6_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_6_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_6_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_6_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_6_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_6_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_7_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_7_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_7_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_7_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_7_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_7_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_7_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_7_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_8_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_8_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_8_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_8_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_8_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_8_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_8_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_8_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_9_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_9_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_9_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_9_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_9_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_9_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_9_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_9_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_10_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_10_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_10_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_10_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_10_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_10_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_10_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_10_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_11_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_11_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_11_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_11_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_11_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_11_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_11_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_11_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_12_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_12_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_12_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_12_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_12_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_12_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_12_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_12_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_13_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_13_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_13_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_13_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_13_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_13_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_13_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_13_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_14_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_14_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_14_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_14_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_14_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_14_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_14_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_14_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_15_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_15_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_15_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_15_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_15_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_15_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_15_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_15_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_in_cnt; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_0; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_1; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_2; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_3; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_4; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_5; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_6; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_7; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_8; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_9; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_10; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_11; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_12; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_13; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_14; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_15; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_clock; // @[PermutationDesigns.scala 48:22]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_in_en; // @[PermutationDesigns.scala 48:22]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_in_cnt; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_0; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_1; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_2; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_3; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_4; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_5; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_6; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_7; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_8; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_9; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_10; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_11; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_12; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_13; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_14; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_15; // @[PermutationDesigns.scala 48:22]
  wire  Permute_switch_w16_bw64_clock; // @[PermutationDesigns.scala 49:24]
  wire  Permute_switch_w16_bw64_reset; // @[PermutationDesigns.scala 49:24]
  wire  Permute_switch_w16_bw64_io_in_valid; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_0; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_1; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_2; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_3; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_4; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_5; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_6; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_7; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_8; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_9; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_10; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_11; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_12; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_13; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_14; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_15; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_0; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_1; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_2; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_3; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_4; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_5; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_6; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_7; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_8; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_9; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_10; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_11; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_12; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_13; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_14; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_15; // @[PermutationDesigns.scala 49:24]
  wire  Permute_switch_w16_bw64_io_in_en; // @[PermutationDesigns.scala 49:24]
  wire  Permute_switch_w16_bw64_io_out_valid; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_0; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_1; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_2; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_3; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_4; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_5; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_6; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_7; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_8; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_9; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_10; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_11; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_12; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_13; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_14; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_15; // @[PermutationDesigns.scala 49:24]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_clock; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_in_en; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_in_cnt; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_0; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_1; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_2; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_3; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_4; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_5; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_6; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_7; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_8; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_9; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_10; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_11; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_12; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_13; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_14; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_15; // @[PermutationDesigns.scala 55:26]
  wire  RAM_Block_N32_w16_bw64_16_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_16_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_16_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_16_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_16_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_16_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_16_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_16_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_17_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_17_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_17_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_17_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_17_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_17_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_17_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_17_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_18_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_18_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_18_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_18_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_18_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_18_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_18_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_18_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_19_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_19_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_19_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_19_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_19_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_19_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_19_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_19_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_20_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_20_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_20_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_20_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_20_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_20_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_20_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_20_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_21_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_21_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_21_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_21_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_21_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_21_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_21_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_21_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_22_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_22_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_22_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_22_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_22_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_22_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_22_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_22_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_23_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_23_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_23_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_23_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_23_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_23_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_23_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_23_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_24_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_24_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_24_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_24_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_24_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_24_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_24_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_24_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_25_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_25_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_25_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_25_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_25_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_25_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_25_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_25_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_26_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_26_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_26_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_26_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_26_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_26_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_26_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_26_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_27_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_27_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_27_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_27_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_27_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_27_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_27_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_27_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_28_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_28_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_28_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_28_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_28_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_28_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_28_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_28_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_29_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_29_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_29_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_29_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_29_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_29_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_29_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_29_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_30_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_30_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_30_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_30_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_30_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_30_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_30_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_30_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_31_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_31_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_31_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_31_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_31_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_31_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_31_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_31_io_out_data; // @[PermutationDesigns.scala 56:41]
  reg [63:0] Perm_shiftregs_data_r; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_1; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_2; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_3; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_4; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_5; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_6; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_7; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_8; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_9; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_10; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_11; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_12; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_13; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_14; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_15; // @[Reg.scala 16:16]
  reg  Perm_shiftregs_valid; // @[Reg.scala 16:16]
  reg  REG; // @[PermutationDesigns.scala 57:47]
  reg  REG_1; // @[PermutationDesigns.scala 57:47]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg [4:0] value_2; // @[Counter.scala 62:40]
  reg [4:0] value_3; // @[Counter.scala 62:40]
  wire  _T_1 = REG & value_2 == 5'h0; // @[PermutationDesigns.scala 61:39]
  reg  r; // @[Reg.scala 16:16]
  wire  _T_3 = REG_1 & value_3 == 5'h0; // @[PermutationDesigns.scala 61:39]
  reg  r_1; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_1; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_2; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_3; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_4; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_5; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_6; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_7; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_8; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_9; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_10; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_11; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_12; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_13; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_14; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_15; // @[Reg.scala 16:16]
  reg  M0_shiftregs_valid; // @[Reg.scala 16:16]
  reg  value_4; // @[Counter.scala 62:40]
  reg  value_5; // @[Counter.scala 62:40]
  reg  value_6; // @[Counter.scala 62:40]
  reg  value_7; // @[Counter.scala 62:40]
  reg  value_9; // @[Counter.scala 62:40]
  reg  PostPC_fullcnt_reg; // @[Reg.scala 16:16]
  reg  PostPC_swtchcnt_reg; // @[Reg.scala 16:16]
  wire  _T_4 = io_in_en & io_in_valid; // @[PermutationDesigns.scala 73:21]
  wire  _value_T_1 = value_4 + 1'h1; // @[Counter.scala 78:24]
  wire  _GEN_39 = value_4 | REG; // @[PermutationDesigns.scala 78:52 80:29 57:47]
  wire  _GEN_47 = io_in_en & io_in_valid ? _GEN_39 : REG; // @[PermutationDesigns.scala 73:35 57:47]
  wire  _value_T_5 = value_5 + 1'h1; // @[Counter.scala 78:24]
  wire  _value_T_9 = value_6 + 1'h1; // @[Counter.scala 78:24]
  wire  _T_19 = io_in_en & Perm_shiftregs_valid; // @[PermutationDesigns.scala 110:21]
  wire  _GEN_63 = PostPC_fullcnt_reg | REG_1; // @[PermutationDesigns.scala 112:54 113:29 57:47]
  wire  _GEN_65 = io_in_en & Perm_shiftregs_valid ? _GEN_63 : REG_1; // @[PermutationDesigns.scala 110:44 57:47]
  wire  wrap_6 = value_2 == 5'h1f; // @[Counter.scala 74:24]
  wire [4:0] _value_T_13 = value_2 + 5'h1; // @[Counter.scala 78:24]
  wire  _value_T_15 = value + 1'h1; // @[Counter.scala 78:24]
  wire  _T_28 = _T_4 & value_4; // @[PermutationDesigns.scala 128:47]
  wire  wrap_8 = value_3 == 5'h1f; // @[Counter.scala 74:24]
  wire [4:0] _value_T_17 = value_3 + 5'h1; // @[Counter.scala 78:24]
  wire  _value_T_19 = value_1 + 1'h1; // @[Counter.scala 78:24]
  wire  _T_37 = _T_19 & PostPC_fullcnt_reg; // @[PermutationDesigns.scala 134:56]
  wire [63:0] _GEN_378 = {{63'd0}, value_4}; // @[PermutationDesigns.scala 161:44]
  wire [64:0] _T_42 = {{1'd0}, _GEN_378}; // @[PermutationDesigns.scala 161:44]
  wire [63:0] _GEN_379 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_0}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_44 = {{1'd0}, _GEN_379}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_380 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_0}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_47 = {{1'd0}, _GEN_380}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_381 = {{63'd0}, value_1}; // @[PermutationDesigns.scala 174:45]
  wire [64:0] _T_49 = {{1'd0}, _GEN_381}; // @[PermutationDesigns.scala 174:45]
  wire [63:0] _GEN_383 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_1}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_53 = {{1'd0}, _GEN_383}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_384 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_1}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_56 = {{1'd0}, _GEN_384}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_387 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_2}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_62 = {{1'd0}, _GEN_387}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_388 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_2}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_65 = {{1'd0}, _GEN_388}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_391 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_3}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_71 = {{1'd0}, _GEN_391}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_392 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_3}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_74 = {{1'd0}, _GEN_392}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_395 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_4}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_80 = {{1'd0}, _GEN_395}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_396 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_4}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_83 = {{1'd0}, _GEN_396}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_399 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_5}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_89 = {{1'd0}, _GEN_399}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_400 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_5}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_92 = {{1'd0}, _GEN_400}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_403 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_6}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_98 = {{1'd0}, _GEN_403}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_404 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_6}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_101 = {{1'd0}, _GEN_404}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_407 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_7}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_107 = {{1'd0}, _GEN_407}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_408 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_7}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_110 = {{1'd0}, _GEN_408}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_411 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_8}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_116 = {{1'd0}, _GEN_411}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_412 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_8}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_119 = {{1'd0}, _GEN_412}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_415 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_9}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_125 = {{1'd0}, _GEN_415}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_416 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_9}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_128 = {{1'd0}, _GEN_416}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_419 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_10}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_134 = {{1'd0}, _GEN_419}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_420 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_10}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_137 = {{1'd0}, _GEN_420}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_423 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_11}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_143 = {{1'd0}, _GEN_423}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_424 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_11}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_146 = {{1'd0}, _GEN_424}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_427 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_12}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_152 = {{1'd0}, _GEN_427}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_428 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_12}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_155 = {{1'd0}, _GEN_428}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_431 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_13}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_161 = {{1'd0}, _GEN_431}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_432 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_13}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_164 = {{1'd0}, _GEN_432}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_435 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_14}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_170 = {{1'd0}, _GEN_435}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_436 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_14}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_173 = {{1'd0}, _GEN_436}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_439 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_15}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_179 = {{1'd0}, _GEN_439}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_440 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_15}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_182 = {{1'd0}, _GEN_440}; // @[PermutationDesigns.scala 173:41]
  reg  out_valid_sr_15; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_240; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_241; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_242; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_243; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_244; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_245; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_246; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_247; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_248; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_249; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_250; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_251; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_252; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_253; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_254; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_255; // @[Reg.scala 16:16]
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_1 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_1_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_1_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_1_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_1_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_1_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_1_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_1_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_1_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_2 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_2_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_2_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_2_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_2_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_2_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_2_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_2_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_2_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_3 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_3_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_3_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_3_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_3_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_3_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_3_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_3_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_3_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_4 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_4_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_4_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_4_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_4_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_4_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_4_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_4_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_4_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_5 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_5_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_5_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_5_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_5_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_5_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_5_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_5_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_5_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_6 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_6_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_6_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_6_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_6_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_6_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_6_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_6_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_6_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_7 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_7_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_7_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_7_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_7_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_7_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_7_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_7_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_7_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_8 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_8_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_8_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_8_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_8_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_8_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_8_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_8_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_8_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_9 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_9_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_9_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_9_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_9_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_9_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_9_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_9_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_9_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_10 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_10_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_10_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_10_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_10_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_10_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_10_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_10_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_10_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_11 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_11_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_11_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_11_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_11_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_11_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_11_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_11_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_11_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_12 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_12_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_12_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_12_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_12_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_12_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_12_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_12_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_12_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_13 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_13_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_13_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_13_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_13_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_13_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_13_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_13_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_13_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_14 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_14_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_14_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_14_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_14_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_14_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_14_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_14_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_14_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_15 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_15_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_15_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_15_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_15_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_15_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_15_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_15_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_15_io_out_data)
  );
  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0 Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0 ( // @[PermutationDesigns.scala 47:25]
    .io_in_cnt(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_in_cnt),
    .io_out_0(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_0),
    .io_out_1(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_1),
    .io_out_2(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_2),
    .io_out_3(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_3),
    .io_out_4(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_4),
    .io_out_5(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_5),
    .io_out_6(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_6),
    .io_out_7(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_7),
    .io_out_8(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_8),
    .io_out_9(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_9),
    .io_out_10(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_10),
    .io_out_11(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_11),
    .io_out_12(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_12),
    .io_out_13(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_13),
    .io_out_14(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_14),
    .io_out_15(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_out_15)
  );
  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1 Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1 ( // @[PermutationDesigns.scala 48:22]
    .clock(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_clock),
    .io_in_en(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_in_en),
    .io_in_cnt(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_in_cnt),
    .io_out_0(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_0),
    .io_out_1(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_1),
    .io_out_2(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_2),
    .io_out_3(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_3),
    .io_out_4(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_4),
    .io_out_5(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_5),
    .io_out_6(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_6),
    .io_out_7(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_7),
    .io_out_8(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_8),
    .io_out_9(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_9),
    .io_out_10(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_10),
    .io_out_11(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_11),
    .io_out_12(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_12),
    .io_out_13(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_13),
    .io_out_14(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_14),
    .io_out_15(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_15)
  );
  Permute_switch_w16_bw64 Permute_switch_w16_bw64 ( // @[PermutationDesigns.scala 49:24]
    .clock(Permute_switch_w16_bw64_clock),
    .reset(Permute_switch_w16_bw64_reset),
    .io_in_valid(Permute_switch_w16_bw64_io_in_valid),
    .io_in_0(Permute_switch_w16_bw64_io_in_0),
    .io_in_1(Permute_switch_w16_bw64_io_in_1),
    .io_in_2(Permute_switch_w16_bw64_io_in_2),
    .io_in_3(Permute_switch_w16_bw64_io_in_3),
    .io_in_4(Permute_switch_w16_bw64_io_in_4),
    .io_in_5(Permute_switch_w16_bw64_io_in_5),
    .io_in_6(Permute_switch_w16_bw64_io_in_6),
    .io_in_7(Permute_switch_w16_bw64_io_in_7),
    .io_in_8(Permute_switch_w16_bw64_io_in_8),
    .io_in_9(Permute_switch_w16_bw64_io_in_9),
    .io_in_10(Permute_switch_w16_bw64_io_in_10),
    .io_in_11(Permute_switch_w16_bw64_io_in_11),
    .io_in_12(Permute_switch_w16_bw64_io_in_12),
    .io_in_13(Permute_switch_w16_bw64_io_in_13),
    .io_in_14(Permute_switch_w16_bw64_io_in_14),
    .io_in_15(Permute_switch_w16_bw64_io_in_15),
    .io_in_config_0(Permute_switch_w16_bw64_io_in_config_0),
    .io_in_config_1(Permute_switch_w16_bw64_io_in_config_1),
    .io_in_config_2(Permute_switch_w16_bw64_io_in_config_2),
    .io_in_config_3(Permute_switch_w16_bw64_io_in_config_3),
    .io_in_config_4(Permute_switch_w16_bw64_io_in_config_4),
    .io_in_config_5(Permute_switch_w16_bw64_io_in_config_5),
    .io_in_config_6(Permute_switch_w16_bw64_io_in_config_6),
    .io_in_config_7(Permute_switch_w16_bw64_io_in_config_7),
    .io_in_config_8(Permute_switch_w16_bw64_io_in_config_8),
    .io_in_config_9(Permute_switch_w16_bw64_io_in_config_9),
    .io_in_config_10(Permute_switch_w16_bw64_io_in_config_10),
    .io_in_config_11(Permute_switch_w16_bw64_io_in_config_11),
    .io_in_config_12(Permute_switch_w16_bw64_io_in_config_12),
    .io_in_config_13(Permute_switch_w16_bw64_io_in_config_13),
    .io_in_config_14(Permute_switch_w16_bw64_io_in_config_14),
    .io_in_config_15(Permute_switch_w16_bw64_io_in_config_15),
    .io_in_en(Permute_switch_w16_bw64_io_in_en),
    .io_out_valid(Permute_switch_w16_bw64_io_out_valid),
    .io_out_0(Permute_switch_w16_bw64_io_out_0),
    .io_out_1(Permute_switch_w16_bw64_io_out_1),
    .io_out_2(Permute_switch_w16_bw64_io_out_2),
    .io_out_3(Permute_switch_w16_bw64_io_out_3),
    .io_out_4(Permute_switch_w16_bw64_io_out_4),
    .io_out_5(Permute_switch_w16_bw64_io_out_5),
    .io_out_6(Permute_switch_w16_bw64_io_out_6),
    .io_out_7(Permute_switch_w16_bw64_io_out_7),
    .io_out_8(Permute_switch_w16_bw64_io_out_8),
    .io_out_9(Permute_switch_w16_bw64_io_out_9),
    .io_out_10(Permute_switch_w16_bw64_io_out_10),
    .io_out_11(Permute_switch_w16_bw64_io_out_11),
    .io_out_12(Permute_switch_w16_bw64_io_out_12),
    .io_out_13(Permute_switch_w16_bw64_io_out_13),
    .io_out_14(Permute_switch_w16_bw64_io_out_14),
    .io_out_15(Permute_switch_w16_bw64_io_out_15)
  );
  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2 Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2 ( // @[PermutationDesigns.scala 55:26]
    .clock(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_clock),
    .io_in_en(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_in_en),
    .io_in_cnt(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_in_cnt),
    .io_out_0(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_0),
    .io_out_1(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_1),
    .io_out_2(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_2),
    .io_out_3(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_3),
    .io_out_4(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_4),
    .io_out_5(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_5),
    .io_out_6(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_6),
    .io_out_7(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_7),
    .io_out_8(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_8),
    .io_out_9(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_9),
    .io_out_10(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_10),
    .io_out_11(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_11),
    .io_out_12(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_12),
    .io_out_13(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_13),
    .io_out_14(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_14),
    .io_out_15(Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_out_15)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_16 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_16_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_16_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_16_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_16_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_16_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_16_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_16_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_16_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_17 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_17_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_17_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_17_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_17_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_17_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_17_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_17_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_17_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_18 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_18_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_18_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_18_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_18_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_18_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_18_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_18_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_18_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_19 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_19_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_19_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_19_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_19_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_19_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_19_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_19_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_19_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_20 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_20_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_20_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_20_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_20_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_20_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_20_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_20_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_20_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_21 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_21_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_21_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_21_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_21_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_21_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_21_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_21_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_21_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_22 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_22_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_22_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_22_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_22_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_22_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_22_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_22_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_22_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_23 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_23_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_23_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_23_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_23_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_23_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_23_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_23_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_23_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_24 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_24_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_24_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_24_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_24_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_24_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_24_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_24_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_24_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_25 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_25_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_25_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_25_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_25_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_25_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_25_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_25_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_25_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_26 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_26_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_26_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_26_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_26_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_26_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_26_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_26_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_26_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_27 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_27_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_27_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_27_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_27_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_27_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_27_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_27_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_27_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_28 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_28_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_28_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_28_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_28_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_28_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_28_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_28_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_28_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_29 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_29_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_29_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_29_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_29_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_29_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_29_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_29_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_29_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_30 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_30_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_30_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_30_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_30_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_30_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_30_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_30_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_30_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_31 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_31_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_31_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_31_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_31_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_31_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_31_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_31_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_31_io_out_data)
  );
  assign io_out_0 = out_data_sr_r_240; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_1 = out_data_sr_r_241; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_2 = out_data_sr_r_242; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_3 = out_data_sr_r_243; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_4 = out_data_sr_r_244; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_5 = out_data_sr_r_245; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_6 = out_data_sr_r_246; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_7 = out_data_sr_r_247; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_8 = out_data_sr_r_248; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_9 = out_data_sr_r_249; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_10 = out_data_sr_r_250; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_11 = out_data_sr_r_251; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_12 = out_data_sr_r_252; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_13 = out_data_sr_r_253; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_14 = out_data_sr_r_254; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_15 = out_data_sr_r_255; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_valid = out_valid_sr_15; // @[PermutationDesigns.scala 182:22]
  assign RAM_Block_N32_w16_bw64_clock = clock;
  assign RAM_Block_N32_w16_bw64_io_in_raddr = _T_44[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_io_in_data = io_in_0; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_1_clock = clock;
  assign RAM_Block_N32_w16_bw64_1_io_in_raddr = _T_53[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_1_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_1_io_in_data = io_in_1; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_1_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_1_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_1_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_2_clock = clock;
  assign RAM_Block_N32_w16_bw64_2_io_in_raddr = _T_62[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_2_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_2_io_in_data = io_in_2; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_2_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_2_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_2_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_3_clock = clock;
  assign RAM_Block_N32_w16_bw64_3_io_in_raddr = _T_71[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_3_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_3_io_in_data = io_in_3; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_3_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_3_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_3_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_4_clock = clock;
  assign RAM_Block_N32_w16_bw64_4_io_in_raddr = _T_80[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_4_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_4_io_in_data = io_in_4; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_4_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_4_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_4_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_5_clock = clock;
  assign RAM_Block_N32_w16_bw64_5_io_in_raddr = _T_89[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_5_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_5_io_in_data = io_in_5; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_5_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_5_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_5_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_6_clock = clock;
  assign RAM_Block_N32_w16_bw64_6_io_in_raddr = _T_98[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_6_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_6_io_in_data = io_in_6; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_6_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_6_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_6_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_7_clock = clock;
  assign RAM_Block_N32_w16_bw64_7_io_in_raddr = _T_107[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_7_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_7_io_in_data = io_in_7; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_7_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_7_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_7_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_8_clock = clock;
  assign RAM_Block_N32_w16_bw64_8_io_in_raddr = _T_116[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_8_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_8_io_in_data = io_in_8; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_8_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_8_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_8_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_9_clock = clock;
  assign RAM_Block_N32_w16_bw64_9_io_in_raddr = _T_125[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_9_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_9_io_in_data = io_in_9; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_9_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_9_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_9_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_10_clock = clock;
  assign RAM_Block_N32_w16_bw64_10_io_in_raddr = _T_134[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_10_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_10_io_in_data = io_in_10; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_10_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_10_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_10_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_11_clock = clock;
  assign RAM_Block_N32_w16_bw64_11_io_in_raddr = _T_143[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_11_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_11_io_in_data = io_in_11; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_11_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_11_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_11_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_12_clock = clock;
  assign RAM_Block_N32_w16_bw64_12_io_in_raddr = _T_152[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_12_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_12_io_in_data = io_in_12; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_12_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_12_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_12_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_13_clock = clock;
  assign RAM_Block_N32_w16_bw64_13_io_in_raddr = _T_161[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_13_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_13_io_in_data = io_in_13; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_13_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_13_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_13_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_14_clock = clock;
  assign RAM_Block_N32_w16_bw64_14_io_in_raddr = _T_170[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_14_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_14_io_in_data = io_in_14; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_14_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_14_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_14_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_15_clock = clock;
  assign RAM_Block_N32_w16_bw64_15_io_in_raddr = _T_179[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_15_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_15_io_in_data = io_in_15; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_15_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_15_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_15_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0_io_in_cnt = value; // @[PermutationDesigns.scala 148:20]
  assign Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_clock = clock;
  assign Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_in_en = io_in_en; // @[PermutationDesigns.scala 150:16]
  assign Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_in_cnt = value_5; // @[PermutationDesigns.scala 152:17]
  assign Permute_switch_w16_bw64_clock = clock;
  assign Permute_switch_w16_bw64_reset = reset;
  assign Permute_switch_w16_bw64_io_in_valid = M0_shiftregs_valid; // @[PermutationDesigns.scala 167:23]
  assign Permute_switch_w16_bw64_io_in_0 = M0_shiftregs_data_r; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_1 = M0_shiftregs_data_r_1; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_2 = M0_shiftregs_data_r_2; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_3 = M0_shiftregs_data_r_3; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_4 = M0_shiftregs_data_r_4; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_5 = M0_shiftregs_data_r_5; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_6 = M0_shiftregs_data_r_6; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_7 = M0_shiftregs_data_r_7; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_8 = M0_shiftregs_data_r_8; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_9 = M0_shiftregs_data_r_9; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_10 = M0_shiftregs_data_r_10; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_11 = M0_shiftregs_data_r_11; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_12 = M0_shiftregs_data_r_12; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_13 = M0_shiftregs_data_r_13; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_14 = M0_shiftregs_data_r_14; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_15 = M0_shiftregs_data_r_15; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_config_0 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_0; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_1 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_1; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_2 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_2; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_3 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_3; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_4 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_4; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_5 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_5; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_6 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_6; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_7 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_7; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_8 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_8; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_9 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_9; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_10 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_10; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_11 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_11; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_12 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_12; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_13 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_13; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_14 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_14; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_15 = Permute_Config_ROM_N32_r2_bitRtrue_w16_stage1_io_out_15; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_en = io_in_en; // @[PermutationDesigns.scala 165:20]
  assign Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_clock = clock;
  assign Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_in_en = io_in_en; // @[PermutationDesigns.scala 153:20]
  assign Permute_Config_ROM_N32_r2_bitRtrue_w16_stage2_io_in_cnt = value_6; // @[PermutationDesigns.scala 155:21]
  assign RAM_Block_N32_w16_bw64_16_clock = clock;
  assign RAM_Block_N32_w16_bw64_16_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_16_io_in_waddr = _T_47[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_16_io_in_data = Perm_shiftregs_data_r; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_16_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_16_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_16_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_17_clock = clock;
  assign RAM_Block_N32_w16_bw64_17_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_17_io_in_waddr = _T_56[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_17_io_in_data = Perm_shiftregs_data_r_1; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_17_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_17_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_17_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_18_clock = clock;
  assign RAM_Block_N32_w16_bw64_18_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_18_io_in_waddr = _T_65[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_18_io_in_data = Perm_shiftregs_data_r_2; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_18_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_18_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_18_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_19_clock = clock;
  assign RAM_Block_N32_w16_bw64_19_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_19_io_in_waddr = _T_74[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_19_io_in_data = Perm_shiftregs_data_r_3; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_19_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_19_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_19_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_20_clock = clock;
  assign RAM_Block_N32_w16_bw64_20_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_20_io_in_waddr = _T_83[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_20_io_in_data = Perm_shiftregs_data_r_4; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_20_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_20_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_20_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_21_clock = clock;
  assign RAM_Block_N32_w16_bw64_21_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_21_io_in_waddr = _T_92[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_21_io_in_data = Perm_shiftregs_data_r_5; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_21_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_21_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_21_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_22_clock = clock;
  assign RAM_Block_N32_w16_bw64_22_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_22_io_in_waddr = _T_101[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_22_io_in_data = Perm_shiftregs_data_r_6; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_22_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_22_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_22_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_23_clock = clock;
  assign RAM_Block_N32_w16_bw64_23_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_23_io_in_waddr = _T_110[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_23_io_in_data = Perm_shiftregs_data_r_7; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_23_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_23_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_23_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_24_clock = clock;
  assign RAM_Block_N32_w16_bw64_24_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_24_io_in_waddr = _T_119[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_24_io_in_data = Perm_shiftregs_data_r_8; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_24_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_24_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_24_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_25_clock = clock;
  assign RAM_Block_N32_w16_bw64_25_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_25_io_in_waddr = _T_128[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_25_io_in_data = Perm_shiftregs_data_r_9; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_25_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_25_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_25_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_26_clock = clock;
  assign RAM_Block_N32_w16_bw64_26_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_26_io_in_waddr = _T_137[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_26_io_in_data = Perm_shiftregs_data_r_10; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_26_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_26_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_26_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_27_clock = clock;
  assign RAM_Block_N32_w16_bw64_27_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_27_io_in_waddr = _T_146[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_27_io_in_data = Perm_shiftregs_data_r_11; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_27_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_27_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_27_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_28_clock = clock;
  assign RAM_Block_N32_w16_bw64_28_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_28_io_in_waddr = _T_155[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_28_io_in_data = Perm_shiftregs_data_r_12; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_28_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_28_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_28_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_29_clock = clock;
  assign RAM_Block_N32_w16_bw64_29_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_29_io_in_waddr = _T_164[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_29_io_in_data = Perm_shiftregs_data_r_13; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_29_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_29_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_29_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_30_clock = clock;
  assign RAM_Block_N32_w16_bw64_30_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_30_io_in_waddr = _T_173[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_30_io_in_data = Perm_shiftregs_data_r_14; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_30_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_30_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_30_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_31_clock = clock;
  assign RAM_Block_N32_w16_bw64_31_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_31_io_in_waddr = _T_182[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_31_io_in_data = Perm_shiftregs_data_r_15; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_31_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_31_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_31_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  always @(posedge clock) begin
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r <= Permute_switch_w16_bw64_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_1 <= Permute_switch_w16_bw64_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_2 <= Permute_switch_w16_bw64_io_out_2; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_3 <= Permute_switch_w16_bw64_io_out_3; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_4 <= Permute_switch_w16_bw64_io_out_4; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_5 <= Permute_switch_w16_bw64_io_out_5; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_6 <= Permute_switch_w16_bw64_io_out_6; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_7 <= Permute_switch_w16_bw64_io_out_7; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_8 <= Permute_switch_w16_bw64_io_out_8; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_9 <= Permute_switch_w16_bw64_io_out_9; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_10 <= Permute_switch_w16_bw64_io_out_10; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_11 <= Permute_switch_w16_bw64_io_out_11; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_12 <= Permute_switch_w16_bw64_io_out_12; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_13 <= Permute_switch_w16_bw64_io_out_13; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_14 <= Permute_switch_w16_bw64_io_out_14; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_15 <= Permute_switch_w16_bw64_io_out_15; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_valid <= Permute_switch_w16_bw64_io_out_valid; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[PermutationDesigns.scala 57:47]
      REG <= 1'h0; // @[PermutationDesigns.scala 57:47]
    end else if (io_in_en & REG) begin // @[PermutationDesigns.scala 119:41]
      if (wrap_6) begin // @[PermutationDesigns.scala 121:57]
        if (value) begin // @[PermutationDesigns.scala 126:57]
          REG <= _T_28;
        end else begin
          REG <= _GEN_47;
        end
      end else begin
        REG <= _GEN_47;
      end
    end else begin
      REG <= _GEN_47;
    end
    if (reset) begin // @[PermutationDesigns.scala 57:47]
      REG_1 <= 1'h0; // @[PermutationDesigns.scala 57:47]
    end else if (io_in_en & REG_1) begin // @[PermutationDesigns.scala 119:41]
      if (wrap_8) begin // @[PermutationDesigns.scala 121:57]
        if (value_1) begin // @[PermutationDesigns.scala 126:57]
          REG_1 <= _T_37;
        end else begin
          REG_1 <= _GEN_65;
        end
      end else begin
        REG_1 <= _GEN_65;
      end
    end else begin
      REG_1 <= _GEN_65;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & REG) begin // @[PermutationDesigns.scala 119:41]
      if (wrap_6) begin // @[PermutationDesigns.scala 121:57]
        value <= _value_T_15;
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & REG_1) begin // @[PermutationDesigns.scala 119:41]
      if (wrap_8) begin // @[PermutationDesigns.scala 121:57]
        value_1 <= _value_T_19;
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_2 <= 5'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & REG) begin // @[PermutationDesigns.scala 119:41]
      value_2 <= _value_T_13; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_3 <= 5'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & REG_1) begin // @[PermutationDesigns.scala 119:41]
      value_3 <= _value_T_17; // @[Counter.scala 78:15]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      r <= _T_1; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      r_1 <= _T_3; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r <= RAM_Block_N32_w16_bw64_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_1 <= RAM_Block_N32_w16_bw64_1_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_2 <= RAM_Block_N32_w16_bw64_2_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_3 <= RAM_Block_N32_w16_bw64_3_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_4 <= RAM_Block_N32_w16_bw64_4_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_5 <= RAM_Block_N32_w16_bw64_5_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_6 <= RAM_Block_N32_w16_bw64_6_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_7 <= RAM_Block_N32_w16_bw64_7_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_8 <= RAM_Block_N32_w16_bw64_8_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_9 <= RAM_Block_N32_w16_bw64_9_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_10 <= RAM_Block_N32_w16_bw64_10_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_11 <= RAM_Block_N32_w16_bw64_11_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_12 <= RAM_Block_N32_w16_bw64_12_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_13 <= RAM_Block_N32_w16_bw64_13_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_14 <= RAM_Block_N32_w16_bw64_14_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_15 <= RAM_Block_N32_w16_bw64_15_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_valid <= r; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_4 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & io_in_valid) begin // @[PermutationDesigns.scala 73:35]
      value_4 <= _value_T_1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_5 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & r) begin // @[PermutationDesigns.scala 86:40]
      value_5 <= _value_T_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_6 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & Permute_switch_w16_bw64_io_out_valid) begin // @[PermutationDesigns.scala 98:38]
      value_6 <= _value_T_9;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_7 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & io_in_valid) begin // @[PermutationDesigns.scala 73:35]
      if (value_4) begin // @[PermutationDesigns.scala 78:52]
        value_7 <= value_7 + 1'h1; // @[Counter.scala 78:15]
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_9 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & Permute_switch_w16_bw64_io_out_valid) begin // @[PermutationDesigns.scala 98:38]
      if (value_6) begin // @[PermutationDesigns.scala 103:52]
        value_9 <= value_9 + 1'h1; // @[Counter.scala 78:15]
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      PostPC_fullcnt_reg <= value_6; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      PostPC_swtchcnt_reg <= value_9; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_valid_sr_15 <= r_1; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_240 <= RAM_Block_N32_w16_bw64_16_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_241 <= RAM_Block_N32_w16_bw64_17_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_242 <= RAM_Block_N32_w16_bw64_18_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_243 <= RAM_Block_N32_w16_bw64_19_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_244 <= RAM_Block_N32_w16_bw64_20_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_245 <= RAM_Block_N32_w16_bw64_21_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_246 <= RAM_Block_N32_w16_bw64_22_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_247 <= RAM_Block_N32_w16_bw64_23_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_248 <= RAM_Block_N32_w16_bw64_24_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_249 <= RAM_Block_N32_w16_bw64_25_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_250 <= RAM_Block_N32_w16_bw64_26_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_251 <= RAM_Block_N32_w16_bw64_27_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_252 <= RAM_Block_N32_w16_bw64_28_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_253 <= RAM_Block_N32_w16_bw64_29_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_254 <= RAM_Block_N32_w16_bw64_30_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_255 <= RAM_Block_N32_w16_bw64_31_io_out_data; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  Perm_shiftregs_data_r = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  Perm_shiftregs_data_r_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  Perm_shiftregs_data_r_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  Perm_shiftregs_data_r_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  Perm_shiftregs_data_r_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  Perm_shiftregs_data_r_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  Perm_shiftregs_data_r_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  Perm_shiftregs_data_r_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  Perm_shiftregs_data_r_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  Perm_shiftregs_data_r_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  Perm_shiftregs_data_r_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  Perm_shiftregs_data_r_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  Perm_shiftregs_data_r_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  Perm_shiftregs_data_r_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  Perm_shiftregs_data_r_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  Perm_shiftregs_data_r_15 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  Perm_shiftregs_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  REG = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  value = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  value_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  value_2 = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  value_3 = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  r = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  r_1 = _RAND_24[0:0];
  _RAND_25 = {2{`RANDOM}};
  M0_shiftregs_data_r = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  M0_shiftregs_data_r_1 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  M0_shiftregs_data_r_2 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  M0_shiftregs_data_r_3 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  M0_shiftregs_data_r_4 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  M0_shiftregs_data_r_5 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  M0_shiftregs_data_r_6 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  M0_shiftregs_data_r_7 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  M0_shiftregs_data_r_8 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  M0_shiftregs_data_r_9 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  M0_shiftregs_data_r_10 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  M0_shiftregs_data_r_11 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  M0_shiftregs_data_r_12 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  M0_shiftregs_data_r_13 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  M0_shiftregs_data_r_14 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  M0_shiftregs_data_r_15 = _RAND_40[63:0];
  _RAND_41 = {1{`RANDOM}};
  M0_shiftregs_valid = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  value_4 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  value_5 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  value_6 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  value_7 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  value_9 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  PostPC_fullcnt_reg = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  PostPC_swtchcnt_reg = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  out_valid_sr_15 = _RAND_49[0:0];
  _RAND_50 = {2{`RANDOM}};
  out_data_sr_r_240 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  out_data_sr_r_241 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  out_data_sr_r_242 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  out_data_sr_r_243 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  out_data_sr_r_244 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  out_data_sr_r_245 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  out_data_sr_r_246 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  out_data_sr_r_247 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  out_data_sr_r_248 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  out_data_sr_r_249 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  out_data_sr_r_250 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  out_data_sr_r_251 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  out_data_sr_r_252 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  out_data_sr_r_253 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  out_data_sr_r_254 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  out_data_sr_r_255 = _RAND_65[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1(
  input        clock,
  input        io_in_en,
  input        io_in_cnt,
  output [3:0] io_out_0,
  output [3:0] io_out_1,
  output [3:0] io_out_2,
  output [3:0] io_out_3,
  output [3:0] io_out_4,
  output [3:0] io_out_5,
  output [3:0] io_out_6,
  output [3:0] io_out_7,
  output [3:0] io_out_8,
  output [3:0] io_out_9,
  output [3:0] io_out_10,
  output [3:0] io_out_11,
  output [3:0] io_out_12,
  output [3:0] io_out_13,
  output [3:0] io_out_14,
  output [3:0] io_out_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] out_reg_data_r; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_1; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_2; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_3; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_4; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_5; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_6; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_7; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_8; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_9; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_10; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_11; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_12; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_13; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_14; // @[Reg.scala 16:16]
  reg [3:0] out_reg_data_r_15; // @[Reg.scala 16:16]
  assign io_out_0 = out_reg_data_r; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_1 = out_reg_data_r_1; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_2 = out_reg_data_r_2; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_3 = out_reg_data_r_3; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_4 = out_reg_data_r_4; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_5 = out_reg_data_r_5; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_6 = out_reg_data_r_6; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_7 = out_reg_data_r_7; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_8 = out_reg_data_r_8; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_9 = out_reg_data_r_9; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_10 = out_reg_data_r_10; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_11 = out_reg_data_r_11; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_12 = out_reg_data_r_12; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_13 = out_reg_data_r_13; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_14 = out_reg_data_r_14; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_15 = out_reg_data_r_15; // @[PermutationDesigns.scala 229:{31,31}]
  always @(posedge clock) begin
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r <= 4'h8; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r <= 4'h0;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_1 <= 4'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_1 <= 4'h8;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_2 <= 4'h9; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_2 <= 4'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_3 <= 4'h1; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_3 <= 4'h9;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_4 <= 4'ha; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_4 <= 4'h2;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_5 <= 4'h2; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_5 <= 4'ha;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_6 <= 4'hb; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_6 <= 4'h3;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_7 <= 4'h3; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_7 <= 4'hb;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_8 <= 4'hc; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_8 <= 4'h4;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_9 <= 4'h4; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_9 <= 4'hc;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_10 <= 4'hd; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_10 <= 4'h5;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_11 <= 4'h5; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_11 <= 4'hd;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_12 <= 4'he; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_12 <= 4'h6;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_13 <= 4'h6; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_13 <= 4'he;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_14 <= 4'hf; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_14 <= 4'h7;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_15 <= 4'h7; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_15 <= 4'hf;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_reg_data_r = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  out_reg_data_r_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  out_reg_data_r_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  out_reg_data_r_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  out_reg_data_r_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  out_reg_data_r_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  out_reg_data_r_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  out_reg_data_r_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  out_reg_data_r_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  out_reg_data_r_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  out_reg_data_r_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  out_reg_data_r_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  out_reg_data_r_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  out_reg_data_r_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  out_reg_data_r_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  out_reg_data_r_15 = _RAND_15[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2(
  input   clock,
  input   io_in_en,
  input   io_in_cnt,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg  out_reg_data_r; // @[Reg.scala 16:16]
  reg  out_reg_data_r_1; // @[Reg.scala 16:16]
  reg  out_reg_data_r_2; // @[Reg.scala 16:16]
  reg  out_reg_data_r_3; // @[Reg.scala 16:16]
  reg  out_reg_data_r_4; // @[Reg.scala 16:16]
  reg  out_reg_data_r_5; // @[Reg.scala 16:16]
  reg  out_reg_data_r_6; // @[Reg.scala 16:16]
  reg  out_reg_data_r_7; // @[Reg.scala 16:16]
  reg  out_reg_data_r_8; // @[Reg.scala 16:16]
  reg  out_reg_data_r_9; // @[Reg.scala 16:16]
  reg  out_reg_data_r_10; // @[Reg.scala 16:16]
  reg  out_reg_data_r_11; // @[Reg.scala 16:16]
  reg  out_reg_data_r_12; // @[Reg.scala 16:16]
  reg  out_reg_data_r_13; // @[Reg.scala 16:16]
  reg  out_reg_data_r_14; // @[Reg.scala 16:16]
  reg  out_reg_data_r_15; // @[Reg.scala 16:16]
  assign io_out_0 = out_reg_data_r; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_1 = out_reg_data_r_1; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_2 = out_reg_data_r_2; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_3 = out_reg_data_r_3; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_4 = out_reg_data_r_4; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_5 = out_reg_data_r_5; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_6 = out_reg_data_r_6; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_7 = out_reg_data_r_7; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_8 = out_reg_data_r_8; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_9 = out_reg_data_r_9; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_10 = out_reg_data_r_10; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_11 = out_reg_data_r_11; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_12 = out_reg_data_r_12; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_13 = out_reg_data_r_13; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_14 = out_reg_data_r_14; // @[PermutationDesigns.scala 229:{31,31}]
  assign io_out_15 = out_reg_data_r_15; // @[PermutationDesigns.scala 229:{31,31}]
  always @(posedge clock) begin
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_1 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_2 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_3 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_4 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_5 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_6 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_reg_data_r_7 <= io_in_cnt; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_8 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_8 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_9 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_9 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_10 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_10 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_11 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_11 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_12 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_12 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_13 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_13 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_14 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_14 <= 1'h1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      if (io_in_cnt) begin // @[Reg.scala 17:22]
        out_reg_data_r_15 <= 1'h0; // @[Reg.scala 17:22]
      end else begin
        out_reg_data_r_15 <= 1'h1;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_reg_data_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_reg_data_r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_reg_data_r_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_reg_data_r_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_reg_data_r_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_reg_data_r_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_reg_data_r_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  out_reg_data_r_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  out_reg_data_r_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  out_reg_data_r_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  out_reg_data_r_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  out_reg_data_r_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  out_reg_data_r_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  out_reg_data_r_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  out_reg_data_r_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  out_reg_data_r_15 = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Permute_Streaming_N32_r2_w16_bitRfalse_bw64(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [63:0] io_in_0,
  input  [63:0] io_in_1,
  input  [63:0] io_in_2,
  input  [63:0] io_in_3,
  input  [63:0] io_in_4,
  input  [63:0] io_in_5,
  input  [63:0] io_in_6,
  input  [63:0] io_in_7,
  input  [63:0] io_in_8,
  input  [63:0] io_in_9,
  input  [63:0] io_in_10,
  input  [63:0] io_in_11,
  input  [63:0] io_in_12,
  input  [63:0] io_in_13,
  input  [63:0] io_in_14,
  input  [63:0] io_in_15,
  input         io_in_valid,
  output [63:0] io_out_0,
  output [63:0] io_out_1,
  output [63:0] io_out_2,
  output [63:0] io_out_3,
  output [63:0] io_out_4,
  output [63:0] io_out_5,
  output [63:0] io_out_6,
  output [63:0] io_out_7,
  output [63:0] io_out_8,
  output [63:0] io_out_9,
  output [63:0] io_out_10,
  output [63:0] io_out_11,
  output [63:0] io_out_12,
  output [63:0] io_out_13,
  output [63:0] io_out_14,
  output [63:0] io_out_15,
  output        io_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_Block_N32_w16_bw64_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_1_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_1_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_1_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_1_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_1_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_1_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_1_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_1_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_2_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_2_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_2_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_2_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_2_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_2_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_2_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_2_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_3_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_3_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_3_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_3_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_3_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_3_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_3_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_3_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_4_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_4_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_4_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_4_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_4_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_4_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_4_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_4_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_5_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_5_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_5_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_5_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_5_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_5_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_5_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_5_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_6_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_6_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_6_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_6_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_6_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_6_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_6_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_6_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_7_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_7_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_7_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_7_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_7_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_7_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_7_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_7_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_8_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_8_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_8_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_8_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_8_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_8_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_8_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_8_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_9_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_9_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_9_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_9_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_9_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_9_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_9_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_9_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_10_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_10_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_10_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_10_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_10_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_10_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_10_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_10_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_11_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_11_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_11_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_11_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_11_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_11_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_11_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_11_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_12_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_12_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_12_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_12_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_12_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_12_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_12_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_12_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_13_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_13_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_13_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_13_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_13_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_13_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_13_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_13_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_14_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_14_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_14_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_14_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_14_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_14_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_14_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_14_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_15_clock; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_15_io_in_raddr; // @[PermutationDesigns.scala 46:37]
  wire [1:0] RAM_Block_N32_w16_bw64_15_io_in_waddr; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_15_io_in_data; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_15_io_in_offset_switch; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_15_io_in_valid; // @[PermutationDesigns.scala 46:37]
  wire  RAM_Block_N32_w16_bw64_15_io_in_en; // @[PermutationDesigns.scala 46:37]
  wire [63:0] RAM_Block_N32_w16_bw64_15_io_out_data; // @[PermutationDesigns.scala 46:37]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_in_cnt; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_0; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_1; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_2; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_3; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_4; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_5; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_6; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_7; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_8; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_9; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_10; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_11; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_12; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_13; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_14; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_15; // @[PermutationDesigns.scala 47:25]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_clock; // @[PermutationDesigns.scala 48:22]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_in_en; // @[PermutationDesigns.scala 48:22]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_in_cnt; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_0; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_1; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_2; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_3; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_4; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_5; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_6; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_7; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_8; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_9; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_10; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_11; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_12; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_13; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_14; // @[PermutationDesigns.scala 48:22]
  wire [3:0] Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_15; // @[PermutationDesigns.scala 48:22]
  wire  Permute_switch_w16_bw64_clock; // @[PermutationDesigns.scala 49:24]
  wire  Permute_switch_w16_bw64_reset; // @[PermutationDesigns.scala 49:24]
  wire  Permute_switch_w16_bw64_io_in_valid; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_0; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_1; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_2; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_3; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_4; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_5; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_6; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_7; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_8; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_9; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_10; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_11; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_12; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_13; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_14; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_in_15; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_0; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_1; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_2; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_3; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_4; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_5; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_6; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_7; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_8; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_9; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_10; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_11; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_12; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_13; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_14; // @[PermutationDesigns.scala 49:24]
  wire [3:0] Permute_switch_w16_bw64_io_in_config_15; // @[PermutationDesigns.scala 49:24]
  wire  Permute_switch_w16_bw64_io_in_en; // @[PermutationDesigns.scala 49:24]
  wire  Permute_switch_w16_bw64_io_out_valid; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_0; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_1; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_2; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_3; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_4; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_5; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_6; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_7; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_8; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_9; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_10; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_11; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_12; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_13; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_14; // @[PermutationDesigns.scala 49:24]
  wire [63:0] Permute_switch_w16_bw64_io_out_15; // @[PermutationDesigns.scala 49:24]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_clock; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_in_en; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_in_cnt; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_0; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_1; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_2; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_3; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_4; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_5; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_6; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_7; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_8; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_9; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_10; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_11; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_12; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_13; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_14; // @[PermutationDesigns.scala 55:26]
  wire  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_15; // @[PermutationDesigns.scala 55:26]
  wire  RAM_Block_N32_w16_bw64_16_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_16_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_16_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_16_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_16_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_16_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_16_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_16_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_17_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_17_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_17_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_17_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_17_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_17_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_17_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_17_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_18_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_18_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_18_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_18_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_18_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_18_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_18_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_18_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_19_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_19_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_19_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_19_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_19_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_19_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_19_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_19_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_20_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_20_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_20_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_20_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_20_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_20_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_20_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_20_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_21_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_21_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_21_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_21_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_21_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_21_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_21_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_21_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_22_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_22_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_22_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_22_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_22_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_22_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_22_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_22_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_23_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_23_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_23_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_23_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_23_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_23_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_23_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_23_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_24_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_24_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_24_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_24_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_24_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_24_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_24_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_24_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_25_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_25_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_25_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_25_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_25_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_25_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_25_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_25_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_26_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_26_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_26_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_26_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_26_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_26_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_26_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_26_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_27_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_27_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_27_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_27_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_27_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_27_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_27_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_27_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_28_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_28_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_28_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_28_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_28_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_28_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_28_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_28_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_29_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_29_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_29_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_29_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_29_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_29_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_29_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_29_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_30_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_30_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_30_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_30_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_30_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_30_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_30_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_30_io_out_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_31_clock; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_31_io_in_raddr; // @[PermutationDesigns.scala 56:41]
  wire [1:0] RAM_Block_N32_w16_bw64_31_io_in_waddr; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_31_io_in_data; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_31_io_in_offset_switch; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_31_io_in_valid; // @[PermutationDesigns.scala 56:41]
  wire  RAM_Block_N32_w16_bw64_31_io_in_en; // @[PermutationDesigns.scala 56:41]
  wire [63:0] RAM_Block_N32_w16_bw64_31_io_out_data; // @[PermutationDesigns.scala 56:41]
  reg [63:0] Perm_shiftregs_data_r; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_1; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_2; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_3; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_4; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_5; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_6; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_7; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_8; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_9; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_10; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_11; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_12; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_13; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_14; // @[Reg.scala 16:16]
  reg [63:0] Perm_shiftregs_data_r_15; // @[Reg.scala 16:16]
  reg  Perm_shiftregs_valid; // @[Reg.scala 16:16]
  reg  REG; // @[PermutationDesigns.scala 57:47]
  reg  REG_1; // @[PermutationDesigns.scala 57:47]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg [4:0] value_2; // @[Counter.scala 62:40]
  reg [4:0] value_3; // @[Counter.scala 62:40]
  wire  _T_1 = REG & value_2 == 5'h0; // @[PermutationDesigns.scala 61:39]
  reg  r; // @[Reg.scala 16:16]
  wire  _T_3 = REG_1 & value_3 == 5'h0; // @[PermutationDesigns.scala 61:39]
  reg  r_1; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_1; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_2; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_3; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_4; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_5; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_6; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_7; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_8; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_9; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_10; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_11; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_12; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_13; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_14; // @[Reg.scala 16:16]
  reg [63:0] M0_shiftregs_data_r_15; // @[Reg.scala 16:16]
  reg  M0_shiftregs_valid; // @[Reg.scala 16:16]
  reg  value_4; // @[Counter.scala 62:40]
  reg  value_5; // @[Counter.scala 62:40]
  reg  value_6; // @[Counter.scala 62:40]
  reg  value_7; // @[Counter.scala 62:40]
  reg  value_9; // @[Counter.scala 62:40]
  reg  PostPC_fullcnt_reg; // @[Reg.scala 16:16]
  reg  PostPC_swtchcnt_reg; // @[Reg.scala 16:16]
  wire  _T_4 = io_in_en & io_in_valid; // @[PermutationDesigns.scala 73:21]
  wire  _value_T_1 = value_4 + 1'h1; // @[Counter.scala 78:24]
  wire  _GEN_39 = value_4 | REG; // @[PermutationDesigns.scala 78:52 80:29 57:47]
  wire  _GEN_47 = io_in_en & io_in_valid ? _GEN_39 : REG; // @[PermutationDesigns.scala 73:35 57:47]
  wire  _value_T_5 = value_5 + 1'h1; // @[Counter.scala 78:24]
  wire  _value_T_9 = value_6 + 1'h1; // @[Counter.scala 78:24]
  wire  _T_19 = io_in_en & Perm_shiftregs_valid; // @[PermutationDesigns.scala 110:21]
  wire  _GEN_63 = PostPC_fullcnt_reg | REG_1; // @[PermutationDesigns.scala 112:54 113:29 57:47]
  wire  _GEN_65 = io_in_en & Perm_shiftregs_valid ? _GEN_63 : REG_1; // @[PermutationDesigns.scala 110:44 57:47]
  wire  wrap_6 = value_2 == 5'h1f; // @[Counter.scala 74:24]
  wire [4:0] _value_T_13 = value_2 + 5'h1; // @[Counter.scala 78:24]
  wire  _value_T_15 = value + 1'h1; // @[Counter.scala 78:24]
  wire  _T_28 = _T_4 & value_4; // @[PermutationDesigns.scala 128:47]
  wire  wrap_8 = value_3 == 5'h1f; // @[Counter.scala 74:24]
  wire [4:0] _value_T_17 = value_3 + 5'h1; // @[Counter.scala 78:24]
  wire  _value_T_19 = value_1 + 1'h1; // @[Counter.scala 78:24]
  wire  _T_37 = _T_19 & PostPC_fullcnt_reg; // @[PermutationDesigns.scala 134:56]
  wire [63:0] _GEN_378 = {{63'd0}, value_4}; // @[PermutationDesigns.scala 161:44]
  wire [64:0] _T_42 = {{1'd0}, _GEN_378}; // @[PermutationDesigns.scala 161:44]
  wire [63:0] _GEN_379 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_0}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_44 = {{1'd0}, _GEN_379}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_380 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_0}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_47 = {{1'd0}, _GEN_380}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_381 = {{63'd0}, value_1}; // @[PermutationDesigns.scala 174:45]
  wire [64:0] _T_49 = {{1'd0}, _GEN_381}; // @[PermutationDesigns.scala 174:45]
  wire [63:0] _GEN_383 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_1}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_53 = {{1'd0}, _GEN_383}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_384 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_1}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_56 = {{1'd0}, _GEN_384}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_387 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_2}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_62 = {{1'd0}, _GEN_387}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_388 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_2}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_65 = {{1'd0}, _GEN_388}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_391 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_3}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_71 = {{1'd0}, _GEN_391}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_392 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_3}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_74 = {{1'd0}, _GEN_392}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_395 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_4}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_80 = {{1'd0}, _GEN_395}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_396 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_4}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_83 = {{1'd0}, _GEN_396}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_399 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_5}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_89 = {{1'd0}, _GEN_399}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_400 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_5}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_92 = {{1'd0}, _GEN_400}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_403 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_6}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_98 = {{1'd0}, _GEN_403}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_404 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_6}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_101 = {{1'd0}, _GEN_404}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_407 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_7}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_107 = {{1'd0}, _GEN_407}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_408 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_7}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_110 = {{1'd0}, _GEN_408}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_411 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_8}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_116 = {{1'd0}, _GEN_411}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_412 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_8}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_119 = {{1'd0}, _GEN_412}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_415 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_9}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_125 = {{1'd0}, _GEN_415}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_416 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_9}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_128 = {{1'd0}, _GEN_416}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_419 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_10}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_134 = {{1'd0}, _GEN_419}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_420 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_10}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_137 = {{1'd0}, _GEN_420}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_423 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_11}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_143 = {{1'd0}, _GEN_423}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_424 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_11}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_146 = {{1'd0}, _GEN_424}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_427 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_12}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_152 = {{1'd0}, _GEN_427}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_428 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_12}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_155 = {{1'd0}, _GEN_428}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_431 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_13}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_161 = {{1'd0}, _GEN_431}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_432 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_13}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_164 = {{1'd0}, _GEN_432}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_435 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_14}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_170 = {{1'd0}, _GEN_435}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_436 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_14}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_173 = {{1'd0}, _GEN_436}; // @[PermutationDesigns.scala 173:41]
  wire [63:0] _GEN_439 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_15}; // @[PermutationDesigns.scala 162:40]
  wire [64:0] _T_179 = {{1'd0}, _GEN_439}; // @[PermutationDesigns.scala 162:40]
  wire [63:0] _GEN_440 = {{63'd0}, Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_15}; // @[PermutationDesigns.scala 173:41]
  wire [64:0] _T_182 = {{1'd0}, _GEN_440}; // @[PermutationDesigns.scala 173:41]
  reg  out_valid_sr_15; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_240; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_241; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_242; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_243; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_244; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_245; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_246; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_247; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_248; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_249; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_250; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_251; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_252; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_253; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_254; // @[Reg.scala 16:16]
  reg [63:0] out_data_sr_r_255; // @[Reg.scala 16:16]
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_1 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_1_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_1_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_1_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_1_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_1_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_1_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_1_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_1_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_2 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_2_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_2_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_2_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_2_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_2_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_2_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_2_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_2_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_3 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_3_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_3_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_3_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_3_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_3_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_3_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_3_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_3_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_4 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_4_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_4_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_4_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_4_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_4_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_4_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_4_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_4_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_5 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_5_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_5_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_5_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_5_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_5_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_5_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_5_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_5_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_6 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_6_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_6_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_6_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_6_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_6_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_6_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_6_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_6_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_7 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_7_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_7_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_7_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_7_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_7_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_7_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_7_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_7_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_8 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_8_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_8_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_8_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_8_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_8_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_8_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_8_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_8_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_9 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_9_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_9_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_9_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_9_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_9_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_9_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_9_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_9_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_10 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_10_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_10_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_10_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_10_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_10_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_10_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_10_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_10_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_11 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_11_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_11_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_11_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_11_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_11_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_11_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_11_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_11_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_12 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_12_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_12_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_12_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_12_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_12_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_12_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_12_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_12_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_13 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_13_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_13_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_13_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_13_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_13_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_13_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_13_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_13_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_14 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_14_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_14_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_14_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_14_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_14_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_14_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_14_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_14_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_15 ( // @[PermutationDesigns.scala 46:37]
    .clock(RAM_Block_N32_w16_bw64_15_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_15_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_15_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_15_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_15_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_15_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_15_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_15_io_out_data)
  );
  Permute_Config_ROM_N32_r2_bitRtrue_w16_stage0 Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0 ( // @[PermutationDesigns.scala 47:25]
    .io_in_cnt(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_in_cnt),
    .io_out_0(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_0),
    .io_out_1(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_1),
    .io_out_2(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_2),
    .io_out_3(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_3),
    .io_out_4(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_4),
    .io_out_5(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_5),
    .io_out_6(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_6),
    .io_out_7(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_7),
    .io_out_8(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_8),
    .io_out_9(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_9),
    .io_out_10(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_10),
    .io_out_11(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_11),
    .io_out_12(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_12),
    .io_out_13(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_13),
    .io_out_14(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_14),
    .io_out_15(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_out_15)
  );
  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1 Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1 ( // @[PermutationDesigns.scala 48:22]
    .clock(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_clock),
    .io_in_en(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_in_en),
    .io_in_cnt(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_in_cnt),
    .io_out_0(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_0),
    .io_out_1(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_1),
    .io_out_2(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_2),
    .io_out_3(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_3),
    .io_out_4(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_4),
    .io_out_5(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_5),
    .io_out_6(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_6),
    .io_out_7(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_7),
    .io_out_8(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_8),
    .io_out_9(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_9),
    .io_out_10(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_10),
    .io_out_11(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_11),
    .io_out_12(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_12),
    .io_out_13(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_13),
    .io_out_14(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_14),
    .io_out_15(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_15)
  );
  Permute_switch_w16_bw64 Permute_switch_w16_bw64 ( // @[PermutationDesigns.scala 49:24]
    .clock(Permute_switch_w16_bw64_clock),
    .reset(Permute_switch_w16_bw64_reset),
    .io_in_valid(Permute_switch_w16_bw64_io_in_valid),
    .io_in_0(Permute_switch_w16_bw64_io_in_0),
    .io_in_1(Permute_switch_w16_bw64_io_in_1),
    .io_in_2(Permute_switch_w16_bw64_io_in_2),
    .io_in_3(Permute_switch_w16_bw64_io_in_3),
    .io_in_4(Permute_switch_w16_bw64_io_in_4),
    .io_in_5(Permute_switch_w16_bw64_io_in_5),
    .io_in_6(Permute_switch_w16_bw64_io_in_6),
    .io_in_7(Permute_switch_w16_bw64_io_in_7),
    .io_in_8(Permute_switch_w16_bw64_io_in_8),
    .io_in_9(Permute_switch_w16_bw64_io_in_9),
    .io_in_10(Permute_switch_w16_bw64_io_in_10),
    .io_in_11(Permute_switch_w16_bw64_io_in_11),
    .io_in_12(Permute_switch_w16_bw64_io_in_12),
    .io_in_13(Permute_switch_w16_bw64_io_in_13),
    .io_in_14(Permute_switch_w16_bw64_io_in_14),
    .io_in_15(Permute_switch_w16_bw64_io_in_15),
    .io_in_config_0(Permute_switch_w16_bw64_io_in_config_0),
    .io_in_config_1(Permute_switch_w16_bw64_io_in_config_1),
    .io_in_config_2(Permute_switch_w16_bw64_io_in_config_2),
    .io_in_config_3(Permute_switch_w16_bw64_io_in_config_3),
    .io_in_config_4(Permute_switch_w16_bw64_io_in_config_4),
    .io_in_config_5(Permute_switch_w16_bw64_io_in_config_5),
    .io_in_config_6(Permute_switch_w16_bw64_io_in_config_6),
    .io_in_config_7(Permute_switch_w16_bw64_io_in_config_7),
    .io_in_config_8(Permute_switch_w16_bw64_io_in_config_8),
    .io_in_config_9(Permute_switch_w16_bw64_io_in_config_9),
    .io_in_config_10(Permute_switch_w16_bw64_io_in_config_10),
    .io_in_config_11(Permute_switch_w16_bw64_io_in_config_11),
    .io_in_config_12(Permute_switch_w16_bw64_io_in_config_12),
    .io_in_config_13(Permute_switch_w16_bw64_io_in_config_13),
    .io_in_config_14(Permute_switch_w16_bw64_io_in_config_14),
    .io_in_config_15(Permute_switch_w16_bw64_io_in_config_15),
    .io_in_en(Permute_switch_w16_bw64_io_in_en),
    .io_out_valid(Permute_switch_w16_bw64_io_out_valid),
    .io_out_0(Permute_switch_w16_bw64_io_out_0),
    .io_out_1(Permute_switch_w16_bw64_io_out_1),
    .io_out_2(Permute_switch_w16_bw64_io_out_2),
    .io_out_3(Permute_switch_w16_bw64_io_out_3),
    .io_out_4(Permute_switch_w16_bw64_io_out_4),
    .io_out_5(Permute_switch_w16_bw64_io_out_5),
    .io_out_6(Permute_switch_w16_bw64_io_out_6),
    .io_out_7(Permute_switch_w16_bw64_io_out_7),
    .io_out_8(Permute_switch_w16_bw64_io_out_8),
    .io_out_9(Permute_switch_w16_bw64_io_out_9),
    .io_out_10(Permute_switch_w16_bw64_io_out_10),
    .io_out_11(Permute_switch_w16_bw64_io_out_11),
    .io_out_12(Permute_switch_w16_bw64_io_out_12),
    .io_out_13(Permute_switch_w16_bw64_io_out_13),
    .io_out_14(Permute_switch_w16_bw64_io_out_14),
    .io_out_15(Permute_switch_w16_bw64_io_out_15)
  );
  Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2 Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2 ( // @[PermutationDesigns.scala 55:26]
    .clock(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_clock),
    .io_in_en(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_in_en),
    .io_in_cnt(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_in_cnt),
    .io_out_0(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_0),
    .io_out_1(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_1),
    .io_out_2(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_2),
    .io_out_3(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_3),
    .io_out_4(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_4),
    .io_out_5(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_5),
    .io_out_6(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_6),
    .io_out_7(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_7),
    .io_out_8(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_8),
    .io_out_9(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_9),
    .io_out_10(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_10),
    .io_out_11(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_11),
    .io_out_12(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_12),
    .io_out_13(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_13),
    .io_out_14(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_14),
    .io_out_15(Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_out_15)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_16 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_16_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_16_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_16_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_16_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_16_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_16_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_16_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_16_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_17 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_17_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_17_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_17_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_17_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_17_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_17_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_17_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_17_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_18 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_18_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_18_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_18_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_18_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_18_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_18_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_18_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_18_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_19 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_19_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_19_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_19_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_19_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_19_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_19_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_19_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_19_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_20 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_20_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_20_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_20_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_20_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_20_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_20_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_20_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_20_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_21 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_21_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_21_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_21_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_21_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_21_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_21_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_21_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_21_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_22 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_22_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_22_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_22_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_22_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_22_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_22_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_22_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_22_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_23 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_23_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_23_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_23_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_23_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_23_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_23_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_23_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_23_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_24 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_24_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_24_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_24_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_24_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_24_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_24_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_24_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_24_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_25 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_25_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_25_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_25_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_25_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_25_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_25_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_25_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_25_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_26 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_26_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_26_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_26_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_26_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_26_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_26_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_26_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_26_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_27 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_27_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_27_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_27_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_27_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_27_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_27_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_27_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_27_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_28 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_28_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_28_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_28_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_28_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_28_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_28_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_28_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_28_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_29 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_29_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_29_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_29_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_29_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_29_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_29_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_29_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_29_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_30 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_30_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_30_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_30_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_30_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_30_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_30_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_30_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_30_io_out_data)
  );
  RAM_Block_N32_w16_bw64 RAM_Block_N32_w16_bw64_31 ( // @[PermutationDesigns.scala 56:41]
    .clock(RAM_Block_N32_w16_bw64_31_clock),
    .io_in_raddr(RAM_Block_N32_w16_bw64_31_io_in_raddr),
    .io_in_waddr(RAM_Block_N32_w16_bw64_31_io_in_waddr),
    .io_in_data(RAM_Block_N32_w16_bw64_31_io_in_data),
    .io_in_offset_switch(RAM_Block_N32_w16_bw64_31_io_in_offset_switch),
    .io_in_valid(RAM_Block_N32_w16_bw64_31_io_in_valid),
    .io_in_en(RAM_Block_N32_w16_bw64_31_io_in_en),
    .io_out_data(RAM_Block_N32_w16_bw64_31_io_out_data)
  );
  assign io_out_0 = out_data_sr_r_240; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_1 = out_data_sr_r_241; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_2 = out_data_sr_r_242; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_3 = out_data_sr_r_243; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_4 = out_data_sr_r_244; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_5 = out_data_sr_r_245; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_6 = out_data_sr_r_246; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_7 = out_data_sr_r_247; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_8 = out_data_sr_r_248; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_9 = out_data_sr_r_249; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_10 = out_data_sr_r_250; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_11 = out_data_sr_r_251; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_12 = out_data_sr_r_252; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_13 = out_data_sr_r_253; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_14 = out_data_sr_r_254; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_15 = out_data_sr_r_255; // @[PermutationDesigns.scala 178:{34,34}]
  assign io_out_valid = out_valid_sr_15; // @[PermutationDesigns.scala 182:22]
  assign RAM_Block_N32_w16_bw64_clock = clock;
  assign RAM_Block_N32_w16_bw64_io_in_raddr = _T_44[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_io_in_data = io_in_0; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_1_clock = clock;
  assign RAM_Block_N32_w16_bw64_1_io_in_raddr = _T_53[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_1_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_1_io_in_data = io_in_1; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_1_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_1_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_1_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_2_clock = clock;
  assign RAM_Block_N32_w16_bw64_2_io_in_raddr = _T_62[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_2_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_2_io_in_data = io_in_2; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_2_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_2_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_2_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_3_clock = clock;
  assign RAM_Block_N32_w16_bw64_3_io_in_raddr = _T_71[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_3_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_3_io_in_data = io_in_3; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_3_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_3_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_3_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_4_clock = clock;
  assign RAM_Block_N32_w16_bw64_4_io_in_raddr = _T_80[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_4_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_4_io_in_data = io_in_4; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_4_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_4_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_4_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_5_clock = clock;
  assign RAM_Block_N32_w16_bw64_5_io_in_raddr = _T_89[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_5_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_5_io_in_data = io_in_5; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_5_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_5_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_5_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_6_clock = clock;
  assign RAM_Block_N32_w16_bw64_6_io_in_raddr = _T_98[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_6_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_6_io_in_data = io_in_6; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_6_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_6_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_6_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_7_clock = clock;
  assign RAM_Block_N32_w16_bw64_7_io_in_raddr = _T_107[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_7_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_7_io_in_data = io_in_7; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_7_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_7_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_7_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_8_clock = clock;
  assign RAM_Block_N32_w16_bw64_8_io_in_raddr = _T_116[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_8_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_8_io_in_data = io_in_8; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_8_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_8_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_8_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_9_clock = clock;
  assign RAM_Block_N32_w16_bw64_9_io_in_raddr = _T_125[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_9_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_9_io_in_data = io_in_9; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_9_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_9_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_9_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_10_clock = clock;
  assign RAM_Block_N32_w16_bw64_10_io_in_raddr = _T_134[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_10_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_10_io_in_data = io_in_10; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_10_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_10_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_10_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_11_clock = clock;
  assign RAM_Block_N32_w16_bw64_11_io_in_raddr = _T_143[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_11_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_11_io_in_data = io_in_11; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_11_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_11_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_11_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_12_clock = clock;
  assign RAM_Block_N32_w16_bw64_12_io_in_raddr = _T_152[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_12_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_12_io_in_data = io_in_12; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_12_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_12_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_12_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_13_clock = clock;
  assign RAM_Block_N32_w16_bw64_13_io_in_raddr = _T_161[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_13_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_13_io_in_data = io_in_13; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_13_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_13_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_13_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_14_clock = clock;
  assign RAM_Block_N32_w16_bw64_14_io_in_raddr = _T_170[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_14_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_14_io_in_data = io_in_14; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_14_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_14_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_14_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign RAM_Block_N32_w16_bw64_15_clock = clock;
  assign RAM_Block_N32_w16_bw64_15_io_in_raddr = _T_179[1:0]; // @[PermutationDesigns.scala 162:24]
  assign RAM_Block_N32_w16_bw64_15_io_in_waddr = _T_42[1:0]; // @[PermutationDesigns.scala 161:24]
  assign RAM_Block_N32_w16_bw64_15_io_in_data = io_in_15; // @[PermutationDesigns.scala 159:23]
  assign RAM_Block_N32_w16_bw64_15_io_in_offset_switch = value_7; // @[PermutationDesigns.scala 163:53]
  assign RAM_Block_N32_w16_bw64_15_io_in_valid = io_in_valid; // @[PermutationDesigns.scala 160:24]
  assign RAM_Block_N32_w16_bw64_15_io_in_en = io_in_en; // @[PermutationDesigns.scala 158:21]
  assign Permute_Config_ROM_N32_r2_bitRfalse_w16_stage0_io_in_cnt = value; // @[PermutationDesigns.scala 148:20]
  assign Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_clock = clock;
  assign Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_in_en = io_in_en; // @[PermutationDesigns.scala 150:16]
  assign Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_in_cnt = value_5; // @[PermutationDesigns.scala 152:17]
  assign Permute_switch_w16_bw64_clock = clock;
  assign Permute_switch_w16_bw64_reset = reset;
  assign Permute_switch_w16_bw64_io_in_valid = M0_shiftregs_valid; // @[PermutationDesigns.scala 167:23]
  assign Permute_switch_w16_bw64_io_in_0 = M0_shiftregs_data_r; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_1 = M0_shiftregs_data_r_1; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_2 = M0_shiftregs_data_r_2; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_3 = M0_shiftregs_data_r_3; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_4 = M0_shiftregs_data_r_4; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_5 = M0_shiftregs_data_r_5; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_6 = M0_shiftregs_data_r_6; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_7 = M0_shiftregs_data_r_7; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_8 = M0_shiftregs_data_r_8; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_9 = M0_shiftregs_data_r_9; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_10 = M0_shiftregs_data_r_10; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_11 = M0_shiftregs_data_r_11; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_12 = M0_shiftregs_data_r_12; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_13 = M0_shiftregs_data_r_13; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_14 = M0_shiftregs_data_r_14; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_15 = M0_shiftregs_data_r_15; // @[PermutationDesigns.scala 63:{38,38}]
  assign Permute_switch_w16_bw64_io_in_config_0 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_0; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_1 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_1; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_2 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_2; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_3 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_3; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_4 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_4; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_5 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_5; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_6 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_6; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_7 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_7; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_8 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_8; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_9 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_9; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_10 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_10; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_11 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_11; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_12 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_12; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_13 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_13; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_14 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_14; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_config_15 = Permute_Config_ROM_N32_r2_bitRfalse_w16_stage1_io_out_15; // @[PermutationDesigns.scala 168:27]
  assign Permute_switch_w16_bw64_io_in_en = io_in_en; // @[PermutationDesigns.scala 165:20]
  assign Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_clock = clock;
  assign Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_in_en = io_in_en; // @[PermutationDesigns.scala 153:20]
  assign Permute_Config_ROM_N32_r2_bitRfalse_w16_stage2_io_in_cnt = value_6; // @[PermutationDesigns.scala 155:21]
  assign RAM_Block_N32_w16_bw64_16_clock = clock;
  assign RAM_Block_N32_w16_bw64_16_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_16_io_in_waddr = _T_47[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_16_io_in_data = Perm_shiftregs_data_r; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_16_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_16_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_16_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_17_clock = clock;
  assign RAM_Block_N32_w16_bw64_17_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_17_io_in_waddr = _T_56[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_17_io_in_data = Perm_shiftregs_data_r_1; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_17_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_17_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_17_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_18_clock = clock;
  assign RAM_Block_N32_w16_bw64_18_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_18_io_in_waddr = _T_65[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_18_io_in_data = Perm_shiftregs_data_r_2; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_18_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_18_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_18_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_19_clock = clock;
  assign RAM_Block_N32_w16_bw64_19_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_19_io_in_waddr = _T_74[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_19_io_in_data = Perm_shiftregs_data_r_3; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_19_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_19_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_19_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_20_clock = clock;
  assign RAM_Block_N32_w16_bw64_20_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_20_io_in_waddr = _T_83[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_20_io_in_data = Perm_shiftregs_data_r_4; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_20_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_20_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_20_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_21_clock = clock;
  assign RAM_Block_N32_w16_bw64_21_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_21_io_in_waddr = _T_92[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_21_io_in_data = Perm_shiftregs_data_r_5; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_21_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_21_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_21_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_22_clock = clock;
  assign RAM_Block_N32_w16_bw64_22_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_22_io_in_waddr = _T_101[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_22_io_in_data = Perm_shiftregs_data_r_6; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_22_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_22_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_22_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_23_clock = clock;
  assign RAM_Block_N32_w16_bw64_23_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_23_io_in_waddr = _T_110[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_23_io_in_data = Perm_shiftregs_data_r_7; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_23_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_23_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_23_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_24_clock = clock;
  assign RAM_Block_N32_w16_bw64_24_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_24_io_in_waddr = _T_119[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_24_io_in_data = Perm_shiftregs_data_r_8; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_24_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_24_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_24_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_25_clock = clock;
  assign RAM_Block_N32_w16_bw64_25_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_25_io_in_waddr = _T_128[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_25_io_in_data = Perm_shiftregs_data_r_9; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_25_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_25_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_25_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_26_clock = clock;
  assign RAM_Block_N32_w16_bw64_26_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_26_io_in_waddr = _T_137[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_26_io_in_data = Perm_shiftregs_data_r_10; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_26_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_26_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_26_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_27_clock = clock;
  assign RAM_Block_N32_w16_bw64_27_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_27_io_in_waddr = _T_146[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_27_io_in_data = Perm_shiftregs_data_r_11; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_27_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_27_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_27_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_28_clock = clock;
  assign RAM_Block_N32_w16_bw64_28_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_28_io_in_waddr = _T_155[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_28_io_in_data = Perm_shiftregs_data_r_12; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_28_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_28_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_28_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_29_clock = clock;
  assign RAM_Block_N32_w16_bw64_29_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_29_io_in_waddr = _T_164[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_29_io_in_data = Perm_shiftregs_data_r_13; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_29_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_29_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_29_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_30_clock = clock;
  assign RAM_Block_N32_w16_bw64_30_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_30_io_in_waddr = _T_173[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_30_io_in_data = Perm_shiftregs_data_r_14; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_30_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_30_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_30_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  assign RAM_Block_N32_w16_bw64_31_clock = clock;
  assign RAM_Block_N32_w16_bw64_31_io_in_raddr = _T_49[1:0]; // @[PermutationDesigns.scala 174:24]
  assign RAM_Block_N32_w16_bw64_31_io_in_waddr = _T_182[1:0]; // @[PermutationDesigns.scala 173:24]
  assign RAM_Block_N32_w16_bw64_31_io_in_data = Perm_shiftregs_data_r_15; // @[PermutationDesigns.scala 50:{40,40}]
  assign RAM_Block_N32_w16_bw64_31_io_in_offset_switch = PostPC_swtchcnt_reg; // @[PermutationDesigns.scala 175:32]
  assign RAM_Block_N32_w16_bw64_31_io_in_valid = Perm_shiftregs_valid; // @[PermutationDesigns.scala 172:24]
  assign RAM_Block_N32_w16_bw64_31_io_in_en = io_in_en; // @[PermutationDesigns.scala 170:21]
  always @(posedge clock) begin
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r <= Permute_switch_w16_bw64_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_1 <= Permute_switch_w16_bw64_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_2 <= Permute_switch_w16_bw64_io_out_2; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_3 <= Permute_switch_w16_bw64_io_out_3; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_4 <= Permute_switch_w16_bw64_io_out_4; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_5 <= Permute_switch_w16_bw64_io_out_5; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_6 <= Permute_switch_w16_bw64_io_out_6; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_7 <= Permute_switch_w16_bw64_io_out_7; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_8 <= Permute_switch_w16_bw64_io_out_8; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_9 <= Permute_switch_w16_bw64_io_out_9; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_10 <= Permute_switch_w16_bw64_io_out_10; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_11 <= Permute_switch_w16_bw64_io_out_11; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_12 <= Permute_switch_w16_bw64_io_out_12; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_13 <= Permute_switch_w16_bw64_io_out_13; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_14 <= Permute_switch_w16_bw64_io_out_14; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_data_r_15 <= Permute_switch_w16_bw64_io_out_15; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      Perm_shiftregs_valid <= Permute_switch_w16_bw64_io_out_valid; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[PermutationDesigns.scala 57:47]
      REG <= 1'h0; // @[PermutationDesigns.scala 57:47]
    end else if (io_in_en & REG) begin // @[PermutationDesigns.scala 119:41]
      if (wrap_6) begin // @[PermutationDesigns.scala 121:57]
        if (value) begin // @[PermutationDesigns.scala 126:57]
          REG <= _T_28;
        end else begin
          REG <= _GEN_47;
        end
      end else begin
        REG <= _GEN_47;
      end
    end else begin
      REG <= _GEN_47;
    end
    if (reset) begin // @[PermutationDesigns.scala 57:47]
      REG_1 <= 1'h0; // @[PermutationDesigns.scala 57:47]
    end else if (io_in_en & REG_1) begin // @[PermutationDesigns.scala 119:41]
      if (wrap_8) begin // @[PermutationDesigns.scala 121:57]
        if (value_1) begin // @[PermutationDesigns.scala 126:57]
          REG_1 <= _T_37;
        end else begin
          REG_1 <= _GEN_65;
        end
      end else begin
        REG_1 <= _GEN_65;
      end
    end else begin
      REG_1 <= _GEN_65;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & REG) begin // @[PermutationDesigns.scala 119:41]
      if (wrap_6) begin // @[PermutationDesigns.scala 121:57]
        value <= _value_T_15;
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & REG_1) begin // @[PermutationDesigns.scala 119:41]
      if (wrap_8) begin // @[PermutationDesigns.scala 121:57]
        value_1 <= _value_T_19;
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_2 <= 5'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & REG) begin // @[PermutationDesigns.scala 119:41]
      value_2 <= _value_T_13; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_3 <= 5'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & REG_1) begin // @[PermutationDesigns.scala 119:41]
      value_3 <= _value_T_17; // @[Counter.scala 78:15]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      r <= _T_1; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      r_1 <= _T_3; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r <= RAM_Block_N32_w16_bw64_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_1 <= RAM_Block_N32_w16_bw64_1_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_2 <= RAM_Block_N32_w16_bw64_2_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_3 <= RAM_Block_N32_w16_bw64_3_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_4 <= RAM_Block_N32_w16_bw64_4_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_5 <= RAM_Block_N32_w16_bw64_5_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_6 <= RAM_Block_N32_w16_bw64_6_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_7 <= RAM_Block_N32_w16_bw64_7_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_8 <= RAM_Block_N32_w16_bw64_8_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_9 <= RAM_Block_N32_w16_bw64_9_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_10 <= RAM_Block_N32_w16_bw64_10_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_11 <= RAM_Block_N32_w16_bw64_11_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_12 <= RAM_Block_N32_w16_bw64_12_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_13 <= RAM_Block_N32_w16_bw64_13_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_14 <= RAM_Block_N32_w16_bw64_14_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_data_r_15 <= RAM_Block_N32_w16_bw64_15_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      M0_shiftregs_valid <= r; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_4 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & io_in_valid) begin // @[PermutationDesigns.scala 73:35]
      value_4 <= _value_T_1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_5 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & r) begin // @[PermutationDesigns.scala 86:40]
      value_5 <= _value_T_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_6 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & Permute_switch_w16_bw64_io_out_valid) begin // @[PermutationDesigns.scala 98:38]
      value_6 <= _value_T_9;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_7 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & io_in_valid) begin // @[PermutationDesigns.scala 73:35]
      if (value_4) begin // @[PermutationDesigns.scala 78:52]
        value_7 <= value_7 + 1'h1; // @[Counter.scala 78:15]
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_9 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en & Permute_switch_w16_bw64_io_out_valid) begin // @[PermutationDesigns.scala 98:38]
      if (value_6) begin // @[PermutationDesigns.scala 103:52]
        value_9 <= value_9 + 1'h1; // @[Counter.scala 78:15]
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      PostPC_fullcnt_reg <= value_6; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      PostPC_swtchcnt_reg <= value_9; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_valid_sr_15 <= r_1; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_240 <= RAM_Block_N32_w16_bw64_16_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_241 <= RAM_Block_N32_w16_bw64_17_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_242 <= RAM_Block_N32_w16_bw64_18_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_243 <= RAM_Block_N32_w16_bw64_19_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_244 <= RAM_Block_N32_w16_bw64_20_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_245 <= RAM_Block_N32_w16_bw64_21_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_246 <= RAM_Block_N32_w16_bw64_22_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_247 <= RAM_Block_N32_w16_bw64_23_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_248 <= RAM_Block_N32_w16_bw64_24_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_249 <= RAM_Block_N32_w16_bw64_25_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_250 <= RAM_Block_N32_w16_bw64_26_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_251 <= RAM_Block_N32_w16_bw64_27_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_252 <= RAM_Block_N32_w16_bw64_28_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_253 <= RAM_Block_N32_w16_bw64_29_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_254 <= RAM_Block_N32_w16_bw64_30_io_out_data; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      out_data_sr_r_255 <= RAM_Block_N32_w16_bw64_31_io_out_data; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  Perm_shiftregs_data_r = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  Perm_shiftregs_data_r_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  Perm_shiftregs_data_r_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  Perm_shiftregs_data_r_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  Perm_shiftregs_data_r_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  Perm_shiftregs_data_r_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  Perm_shiftregs_data_r_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  Perm_shiftregs_data_r_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  Perm_shiftregs_data_r_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  Perm_shiftregs_data_r_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  Perm_shiftregs_data_r_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  Perm_shiftregs_data_r_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  Perm_shiftregs_data_r_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  Perm_shiftregs_data_r_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  Perm_shiftregs_data_r_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  Perm_shiftregs_data_r_15 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  Perm_shiftregs_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  REG = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  value = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  value_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  value_2 = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  value_3 = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  r = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  r_1 = _RAND_24[0:0];
  _RAND_25 = {2{`RANDOM}};
  M0_shiftregs_data_r = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  M0_shiftregs_data_r_1 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  M0_shiftregs_data_r_2 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  M0_shiftregs_data_r_3 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  M0_shiftregs_data_r_4 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  M0_shiftregs_data_r_5 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  M0_shiftregs_data_r_6 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  M0_shiftregs_data_r_7 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  M0_shiftregs_data_r_8 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  M0_shiftregs_data_r_9 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  M0_shiftregs_data_r_10 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  M0_shiftregs_data_r_11 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  M0_shiftregs_data_r_12 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  M0_shiftregs_data_r_13 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  M0_shiftregs_data_r_14 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  M0_shiftregs_data_r_15 = _RAND_40[63:0];
  _RAND_41 = {1{`RANDOM}};
  M0_shiftregs_valid = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  value_4 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  value_5 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  value_6 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  value_7 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  value_9 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  PostPC_fullcnt_reg = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  PostPC_swtchcnt_reg = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  out_valid_sr_15 = _RAND_49[0:0];
  _RAND_50 = {2{`RANDOM}};
  out_data_sr_r_240 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  out_data_sr_r_241 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  out_data_sr_r_242 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  out_data_sr_r_243 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  out_data_sr_r_244 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  out_data_sr_r_245 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  out_data_sr_r_246 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  out_data_sr_r_247 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  out_data_sr_r_248 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  out_data_sr_r_249 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  out_data_sr_r_250 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  out_data_sr_r_251 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  out_data_sr_r_252 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  out_data_sr_r_253 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  out_data_sr_r_254 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  out_data_sr_r_255 = _RAND_65[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32(
  input         io_in_inv,
  input  [4:0]  io_in_addr,
  output [31:0] io_out_data_0_Im,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_2_Im,
  output [31:0] io_out_data_3_Re,
  output [31:0] io_out_data_3_Im,
  output [31:0] io_out_data_4_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_6_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im,
  output [31:0] io_out_data_8_Im,
  output [31:0] io_out_data_9_Re,
  output [31:0] io_out_data_9_Im,
  output [31:0] io_out_data_10_Im,
  output [31:0] io_out_data_11_Re,
  output [31:0] io_out_data_11_Im,
  output [31:0] io_out_data_12_Im,
  output [31:0] io_out_data_13_Re,
  output [31:0] io_out_data_13_Im,
  output [31:0] io_out_data_14_Im,
  output [31:0] io_out_data_15_Re,
  output [31:0] io_out_data_15_Im
);
  wire [31:0] _GEN_10 = io_in_addr[0] ? 32'hbe14fdf0 : 32'h3f800000; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_11 = io_in_addr[0] ? 32'h3f7d4694 : 32'h0; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_14 = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_15 = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[TwidFactorDesigns.scala 26:{53,53}]
  assign io_out_data_0_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_1_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_1_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_2_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_3_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_3_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_4_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_5_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_5_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_6_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_7_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_7_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_8_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_9_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_9_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_10_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_11_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_11_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_12_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_13_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_13_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_14_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_15_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_15_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
endmodule
module ComplexMULT_SCAL_NOFP_bw32(
  input  [31:0] io_in_Re,
  input  [31:0] io_in_Im,
  input         io_in_en,
  input         io_is_neg,
  input         io_is_flip,
  output [31:0] io_out_Re,
  output [31:0] io_out_Im
);
  wire  sign_0 = io_in_Re[31]; // @[FPComplex.scala 434:24]
  wire  sign_1 = io_in_Im[31]; // @[FPComplex.scala 435:24]
  wire [7:0] exp_0 = io_in_Re[30:23]; // @[FPComplex.scala 437:23]
  wire [7:0] exp_1 = io_in_Im[30:23]; // @[FPComplex.scala 438:23]
  wire [22:0] frac_0 = io_in_Re[22:0]; // @[FPComplex.scala 440:24]
  wire [22:0] frac_1 = io_in_Im[22:0]; // @[FPComplex.scala 441:24]
  wire  new_sign_0 = io_is_neg ? ~sign_0 : sign_0; // @[FPComplex.scala 443:21 444:19 447:19]
  wire  new_sign_1 = io_is_neg ? ~sign_1 : sign_1; // @[FPComplex.scala 443:21 445:19 448:19]
  wire [7:0] _new_exp_0_T_1 = exp_0 - 8'h0; // @[FPComplex.scala 452:28]
  wire [7:0] new_exp_0 = exp_0 != 8'h0 ? _new_exp_0_T_1 : exp_0; // @[FPComplex.scala 451:26 452:18 454:18]
  wire [7:0] _new_exp_1_T_1 = exp_1 - 8'h0; // @[FPComplex.scala 457:28]
  wire [7:0] new_exp_1 = exp_1 != 8'h0 ? _new_exp_1_T_1 : exp_1; // @[FPComplex.scala 456:26 457:18 459:18]
  wire  _io_out_Re_T = ~new_sign_1; // @[FPComplex.scala 465:23]
  wire [31:0] _io_out_Re_T_2 = {_io_out_Re_T,new_exp_1,frac_1}; // @[FPComplex.scala 465:51]
  wire [31:0] _io_out_Im_T_1 = {new_sign_0,new_exp_0,frac_0}; // @[FPComplex.scala 466:48]
  wire [31:0] _io_out_Im_T_3 = {new_sign_1,new_exp_1,frac_1}; // @[FPComplex.scala 469:48]
  wire [31:0] _GEN_4 = io_is_flip ? _io_out_Re_T_2 : _io_out_Im_T_1; // @[FPComplex.scala 464:23 465:19 468:19]
  wire [31:0] _GEN_5 = io_is_flip ? _io_out_Im_T_1 : _io_out_Im_T_3; // @[FPComplex.scala 464:23 466:19 469:19]
  assign io_out_Re = io_in_en ? _GEN_4 : 32'h0; // @[FPComplex.scala 461:15 463:19]
  assign io_out_Im = io_in_en ? _GEN_5 : 32'h0; // @[FPComplex.scala 462:15 463:19]
endmodule
module TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32(
  input         clock,
  input         reset,
  input         io_in_inv,
  input         io_in_en,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_valid,
  output        io_out_valid,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
`endif // RANDOMIZE_REG_INIT
  wire  TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_inv; // @[TwidFactorDesigns.scala 49:28]
  wire [4:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_addr; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_0_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_1_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_1_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_2_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_3_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_3_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_4_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_5_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_5_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_6_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_7_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_7_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_8_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_9_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_9_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_10_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_11_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_11_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_12_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_13_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_13_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_14_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_15_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_15_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_1_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_1_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_1_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_1_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_1_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_1_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_1_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_2_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_2_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_2_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_2_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_2_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_2_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_2_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_3_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_3_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_3_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_3_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_3_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_3_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_3_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_4_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_4_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_4_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_4_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_4_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_4_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_4_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_5_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_5_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_5_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_5_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_5_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_5_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_5_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_6_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_6_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_6_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_6_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_6_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_6_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_6_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_7_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_7_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_7_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_7_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_7_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_7_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_7_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_8_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_8_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_8_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_8_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_8_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_8_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_8_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_9_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_9_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_9_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_9_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_9_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_9_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_9_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_10_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_10_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_10_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_10_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_10_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_10_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_10_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_11_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_11_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_11_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_11_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_11_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_11_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_11_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_12_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_12_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_12_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_12_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_12_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_12_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_12_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_13_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_13_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_13_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_13_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_13_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_13_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_13_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_14_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_14_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_14_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_14_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_14_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_14_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_14_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_15_io_in_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_15_io_in_Im; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_15_io_in_en; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_15_io_is_neg; // @[TwidFactorDesigns.scala 81:32]
  wire  ComplexMULT_SCAL_NOFP_bw32_15_io_is_flip; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_15_io_out_Re; // @[TwidFactorDesigns.scala 81:32]
  wire [31:0] ComplexMULT_SCAL_NOFP_bw32_15_io_out_Im; // @[TwidFactorDesigns.scala 81:32]
  reg  value_1; // @[Counter.scala 62:40]
  wire  _value_T_1 = value_1 + 1'h1; // @[Counter.scala 78:24]
  wire [63:0] _T_1 = {32'h3f800000,TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_0_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_16 = {TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_1_Re,
    TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_1_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_31 = {32'h3f800000,TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_2_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_46 = {TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_3_Re,
    TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_3_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_61 = {32'h3f800000,TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_4_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_76 = {TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_5_Re,
    TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_5_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_91 = {32'h3f800000,TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_6_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_106 = {TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_7_Re,
    TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_7_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_121 = {32'h3f800000,TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_8_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_136 = {TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_9_Re,
    TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_9_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_151 = {32'h3f800000,TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_10_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_166 = {TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_11_Re,
    TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_11_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_181 = {32'h3f800000,TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_12_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_196 = {TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_13_Re,
    TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_13_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_211 = {32'h3f800000,TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_14_Im}; // @[TwidFactorDesigns.scala 88:45]
  wire [63:0] _T_226 = {TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_15_Re,
    TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_15_Im}; // @[TwidFactorDesigns.scala 88:45]
  reg [31:0] sr_result_regs_r_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_1_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_1_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_2_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_2_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_3_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_3_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_4_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_4_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_5_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_5_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_6_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_6_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_7_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_7_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_8_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_8_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_9_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_9_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_10_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_10_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_11_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_11_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_12_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_12_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_13_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_13_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_14_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_14_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_15_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_15_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_16_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_16_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_17_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_17_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_18_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_18_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_19_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_19_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_20_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_20_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_21_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_21_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_22_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_22_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_23_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_23_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_24_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_24_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_25_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_25_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_26_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_26_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_27_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_27_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_28_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_28_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_29_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_29_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_30_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_30_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_31_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_31_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_32_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_32_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_33_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_33_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_34_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_34_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_35_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_35_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_36_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_36_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_37_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_37_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_38_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_38_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_39_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_39_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_40_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_40_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_41_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_41_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_42_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_42_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_43_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_43_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_44_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_44_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_45_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_45_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_46_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_46_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_47_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_47_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_48_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_48_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_49_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_49_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_50_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_50_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_51_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_51_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_52_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_52_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_53_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_53_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_54_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_54_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_55_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_55_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_56_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_56_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_57_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_57_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_58_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_58_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_59_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_59_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_60_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_60_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_61_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_61_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_62_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_62_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_63_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_63_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_64_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_64_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_65_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_65_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_66_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_66_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_67_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_67_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_68_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_68_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_69_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_69_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_70_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_70_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_71_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_71_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_72_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_72_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_73_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_73_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_74_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_74_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_75_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_75_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_76_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_76_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_77_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_77_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_78_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_78_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_79_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_79_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_80_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_80_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_81_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_81_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_82_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_82_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_83_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_83_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_84_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_84_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_85_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_85_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_86_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_86_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_87_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_87_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_88_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_88_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_89_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_89_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_90_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_90_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_91_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_91_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_92_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_92_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_93_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_93_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_94_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_94_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_95_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_95_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_96_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_96_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_97_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_97_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_98_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_98_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_99_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_99_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_100_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_100_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_101_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_101_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_102_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_102_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_103_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_103_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_104_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_104_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_105_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_105_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_106_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_106_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_107_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_107_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_108_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_108_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_109_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_109_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_110_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_110_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_111_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_111_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_112_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_112_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_113_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_113_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_114_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_114_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_115_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_115_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_116_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_116_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_117_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_117_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_118_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_118_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_119_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_119_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_120_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_120_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_121_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_121_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_122_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_122_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_123_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_123_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_124_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_124_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_125_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_125_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_126_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_126_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_127_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_127_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_128_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_128_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_129_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_129_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_130_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_130_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_131_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_131_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_132_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_132_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_133_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_133_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_134_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_134_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_135_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_135_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_136_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_136_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_137_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_137_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_138_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_138_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_139_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_139_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_140_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_140_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_141_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_141_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_142_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_142_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_143_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_143_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_144_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_144_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_145_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_145_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_146_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_146_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_147_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_147_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_148_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_148_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_149_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_149_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_150_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_150_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_151_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_151_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_152_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_152_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_153_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_153_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_154_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_154_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_155_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_155_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_156_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_156_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_157_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_157_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_158_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_158_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_159_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_159_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_160_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_160_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_161_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_161_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_162_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_162_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_163_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_163_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_164_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_164_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_165_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_165_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_166_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_166_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_167_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_167_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_168_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_168_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_169_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_169_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_170_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_170_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_171_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_171_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_172_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_172_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_173_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_173_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_174_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_174_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_175_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_175_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_176_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_176_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_177_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_177_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_178_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_178_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_179_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_179_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_180_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_180_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_181_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_181_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_182_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_182_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_183_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_183_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_184_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_184_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_185_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_185_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_186_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_186_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_187_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_187_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_188_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_188_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_189_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_189_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_190_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_190_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_191_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_191_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_192_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_192_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_193_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_193_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_194_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_194_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_195_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_195_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_196_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_196_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_197_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_197_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_198_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_198_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_199_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_199_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_200_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_200_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_201_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_201_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_202_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_202_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_203_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_203_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_204_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_204_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_205_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_205_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_206_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_206_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_207_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_207_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_208_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_208_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_209_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_209_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_210_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_210_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_211_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_211_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_212_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_212_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_213_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_213_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_214_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_214_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_215_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_215_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_216_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_216_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_217_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_217_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_218_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_218_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_219_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_219_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_220_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_220_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_221_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_221_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_222_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_222_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_223_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_223_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_224_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_224_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_225_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_225_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_226_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_226_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_227_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_227_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_228_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_228_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_229_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_229_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_230_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_230_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_231_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_231_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_232_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_232_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_233_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_233_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_234_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_234_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_235_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_235_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_236_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_236_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_237_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_237_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_238_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_238_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_239_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_239_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_240_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_240_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_241_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_241_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_242_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_242_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_243_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_243_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_244_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_244_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_245_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_245_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_246_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_246_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_247_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_247_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_248_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_248_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_249_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_249_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_250_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_250_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_251_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_251_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_252_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_252_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_253_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_253_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_254_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_254_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_255_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_255_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_256_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_256_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_257_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_257_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_258_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_258_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_259_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_259_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_260_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_260_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_261_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_261_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_262_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_262_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_263_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_263_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_264_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_264_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_265_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_265_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_266_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_266_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_267_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_267_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_268_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_268_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_269_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_269_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_270_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_270_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_271_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_271_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_272_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_272_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_273_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_273_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_274_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_274_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_275_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_275_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_276_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_276_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_277_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_277_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_278_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_278_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_279_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_279_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_280_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_280_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_281_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_281_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_282_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_282_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_283_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_283_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_284_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_284_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_285_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_285_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_286_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_286_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_287_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_287_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_288_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_288_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_289_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_289_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_290_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_290_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_291_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_291_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_292_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_292_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_293_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_293_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_294_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_294_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_295_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_295_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_296_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_296_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_297_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_297_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_298_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_298_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_299_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_299_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_300_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_300_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_301_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_301_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_302_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_302_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_303_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_303_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_304_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_304_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_305_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_305_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_306_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_306_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_307_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_307_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_308_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_308_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_309_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_309_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_310_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_310_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_311_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_311_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_312_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_312_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_313_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_313_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_314_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_314_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_315_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_315_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_316_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_316_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_317_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_317_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_318_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_318_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_319_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_319_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_320_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_320_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_321_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_321_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_322_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_322_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_323_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_323_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_324_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_324_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_325_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_325_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_326_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_326_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_327_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_327_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_328_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_328_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_329_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_329_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_330_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_330_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_331_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_331_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_332_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_332_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_333_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_333_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_334_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_334_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_335_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_335_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_336_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_336_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_337_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_337_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_338_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_338_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_339_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_339_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_340_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_340_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_341_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_341_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_342_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_342_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_343_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_343_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_344_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_344_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_345_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_345_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_346_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_346_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_347_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_347_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_348_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_348_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_349_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_349_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_350_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_350_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_351_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_351_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_352_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_352_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_353_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_353_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_354_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_354_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_355_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_355_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_356_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_356_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_357_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_357_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_358_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_358_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_359_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_359_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_360_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_360_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_361_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_361_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_362_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_362_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_363_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_363_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_364_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_364_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_365_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_365_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_366_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_366_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_367_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_367_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_368_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_368_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_369_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_369_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_370_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_370_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_371_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_371_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_372_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_372_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_373_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_373_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_374_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_374_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_375_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_375_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_376_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_376_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_377_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_377_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_378_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_378_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_379_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_379_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_380_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_380_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_381_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_381_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_382_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_382_Im; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_383_Re; // @[Reg.scala 16:16]
  reg [31:0] sr_result_regs_r_383_Im; // @[Reg.scala 16:16]
  reg  io_out_valid_r; // @[Reg.scala 16:16]
  reg  io_out_valid_r_1; // @[Reg.scala 16:16]
  reg  io_out_valid_r_2; // @[Reg.scala 16:16]
  reg  io_out_valid_r_3; // @[Reg.scala 16:16]
  reg  io_out_valid_r_4; // @[Reg.scala 16:16]
  reg  io_out_valid_r_5; // @[Reg.scala 16:16]
  reg  io_out_valid_r_6; // @[Reg.scala 16:16]
  reg  io_out_valid_r_7; // @[Reg.scala 16:16]
  reg  io_out_valid_r_8; // @[Reg.scala 16:16]
  reg  io_out_valid_r_9; // @[Reg.scala 16:16]
  reg  io_out_valid_r_10; // @[Reg.scala 16:16]
  reg  io_out_valid_r_11; // @[Reg.scala 16:16]
  reg  io_out_valid_r_12; // @[Reg.scala 16:16]
  reg  io_out_valid_r_13; // @[Reg.scala 16:16]
  reg  io_out_valid_r_14; // @[Reg.scala 16:16]
  reg  io_out_valid_r_15; // @[Reg.scala 16:16]
  reg  io_out_valid_r_16; // @[Reg.scala 16:16]
  reg  io_out_valid_r_17; // @[Reg.scala 16:16]
  reg  io_out_valid_r_18; // @[Reg.scala 16:16]
  reg  io_out_valid_r_19; // @[Reg.scala 16:16]
  reg  io_out_valid_r_20; // @[Reg.scala 16:16]
  reg  io_out_valid_r_21; // @[Reg.scala 16:16]
  reg  io_out_valid_r_22; // @[Reg.scala 16:16]
  reg  io_out_valid_r_23; // @[Reg.scala 16:16]
  TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32 TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32 ( // @[TwidFactorDesigns.scala 49:28]
    .io_in_inv(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_inv),
    .io_in_addr(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_addr),
    .io_out_data_0_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_0_Im),
    .io_out_data_1_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_1_Im),
    .io_out_data_2_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_2_Im),
    .io_out_data_3_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_3_Re),
    .io_out_data_3_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_3_Im),
    .io_out_data_4_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_4_Im),
    .io_out_data_5_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_5_Im),
    .io_out_data_6_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_6_Im),
    .io_out_data_7_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_7_Im),
    .io_out_data_8_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_8_Im),
    .io_out_data_9_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_9_Re),
    .io_out_data_9_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_9_Im),
    .io_out_data_10_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_10_Im),
    .io_out_data_11_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_11_Re),
    .io_out_data_11_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_11_Im),
    .io_out_data_12_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_12_Im),
    .io_out_data_13_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_13_Re),
    .io_out_data_13_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_13_Im),
    .io_out_data_14_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_14_Im),
    .io_out_data_15_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_15_Re),
    .io_out_data_15_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_data_15_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_1 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_1_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_1_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_1_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_1_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_1_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_1_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_1_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_2 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_2_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_2_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_2_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_2_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_2_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_2_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_2_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_3 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_3_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_3_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_3_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_3_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_3_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_3_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_3_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_4 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_4_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_4_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_4_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_4_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_4_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_4_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_4_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_5 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_5_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_5_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_5_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_5_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_5_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_5_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_5_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_6 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_6_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_6_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_6_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_6_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_6_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_6_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_6_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_7 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_7_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_7_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_7_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_7_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_7_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_7_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_7_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_8 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_8_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_8_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_8_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_8_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_8_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_8_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_8_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_9 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_9_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_9_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_9_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_9_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_9_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_9_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_9_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_10 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_10_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_10_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_10_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_10_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_10_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_10_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_10_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_11 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_11_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_11_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_11_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_11_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_11_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_11_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_11_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_12 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_12_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_12_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_12_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_12_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_12_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_12_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_12_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_13 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_13_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_13_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_13_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_13_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_13_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_13_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_13_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_14 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_14_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_14_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_14_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_14_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_14_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_14_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_14_io_out_Im)
  );
  ComplexMULT_SCAL_NOFP_bw32 ComplexMULT_SCAL_NOFP_bw32_15 ( // @[TwidFactorDesigns.scala 81:32]
    .io_in_Re(ComplexMULT_SCAL_NOFP_bw32_15_io_in_Re),
    .io_in_Im(ComplexMULT_SCAL_NOFP_bw32_15_io_in_Im),
    .io_in_en(ComplexMULT_SCAL_NOFP_bw32_15_io_in_en),
    .io_is_neg(ComplexMULT_SCAL_NOFP_bw32_15_io_is_neg),
    .io_is_flip(ComplexMULT_SCAL_NOFP_bw32_15_io_is_flip),
    .io_out_Re(ComplexMULT_SCAL_NOFP_bw32_15_io_out_Re),
    .io_out_Im(ComplexMULT_SCAL_NOFP_bw32_15_io_out_Im)
  );
  assign io_out_valid = io_out_valid_r_23; // @[TwidFactorDesigns.scala 108:22]
  assign io_out_0_Re = sr_result_regs_r_23_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_0_Im = sr_result_regs_r_23_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_1_Re = sr_result_regs_r_47_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_1_Im = sr_result_regs_r_47_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_2_Re = sr_result_regs_r_71_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_2_Im = sr_result_regs_r_71_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_3_Re = sr_result_regs_r_95_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_3_Im = sr_result_regs_r_95_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_4_Re = sr_result_regs_r_119_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_4_Im = sr_result_regs_r_119_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_5_Re = sr_result_regs_r_143_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_5_Im = sr_result_regs_r_143_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_6_Re = sr_result_regs_r_167_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_6_Im = sr_result_regs_r_167_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_7_Re = sr_result_regs_r_191_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_7_Im = sr_result_regs_r_191_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_8_Re = sr_result_regs_r_215_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_8_Im = sr_result_regs_r_215_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_9_Re = sr_result_regs_r_239_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_9_Im = sr_result_regs_r_239_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_10_Re = sr_result_regs_r_263_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_10_Im = sr_result_regs_r_263_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_11_Re = sr_result_regs_r_287_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_11_Im = sr_result_regs_r_287_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_12_Re = sr_result_regs_r_311_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_12_Im = sr_result_regs_r_311_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_13_Re = sr_result_regs_r_335_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_13_Im = sr_result_regs_r_335_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_14_Re = sr_result_regs_r_359_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_14_Im = sr_result_regs_r_359_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_15_Re = sr_result_regs_r_383_Re; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign io_out_15_Im = sr_result_regs_r_383_Im; // @[TwidFactorDesigns.scala 104:{37,37}]
  assign TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_inv = io_in_inv; // @[TwidFactorDesigns.scala 56:23]
  assign TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_addr = {{4'd0}, value_1}; // @[TwidFactorDesigns.scala 55:24]
  assign ComplexMULT_SCAL_NOFP_bw32_io_in_Re = io_in_0_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_io_in_Im = io_in_0_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_io_is_neg = _T_1[62:32] == 31'h3f800000 ? _T_1[63] : _T_1[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_io_is_flip = _T_1[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_1_io_in_Re = io_in_1_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_1_io_in_Im = io_in_1_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_1_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_1_io_is_neg = _T_16[62:32] == 31'h3f800000 ? _T_16[63] : _T_16[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_1_io_is_flip = _T_16[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_2_io_in_Re = io_in_2_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_2_io_in_Im = io_in_2_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_2_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_2_io_is_neg = _T_31[62:32] == 31'h3f800000 ? _T_31[63] : _T_31[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_2_io_is_flip = _T_31[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_3_io_in_Re = io_in_3_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_3_io_in_Im = io_in_3_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_3_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_3_io_is_neg = _T_46[62:32] == 31'h3f800000 ? _T_46[63] : _T_46[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_3_io_is_flip = _T_46[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_4_io_in_Re = io_in_4_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_4_io_in_Im = io_in_4_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_4_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_4_io_is_neg = _T_61[62:32] == 31'h3f800000 ? _T_61[63] : _T_61[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_4_io_is_flip = _T_61[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_5_io_in_Re = io_in_5_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_5_io_in_Im = io_in_5_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_5_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_5_io_is_neg = _T_76[62:32] == 31'h3f800000 ? _T_76[63] : _T_76[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_5_io_is_flip = _T_76[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_6_io_in_Re = io_in_6_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_6_io_in_Im = io_in_6_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_6_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_6_io_is_neg = _T_91[62:32] == 31'h3f800000 ? _T_91[63] : _T_91[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_6_io_is_flip = _T_91[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_7_io_in_Re = io_in_7_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_7_io_in_Im = io_in_7_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_7_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_7_io_is_neg = _T_106[62:32] == 31'h3f800000 ? _T_106[63] : _T_106[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_7_io_is_flip = _T_106[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_8_io_in_Re = io_in_8_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_8_io_in_Im = io_in_8_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_8_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_8_io_is_neg = _T_121[62:32] == 31'h3f800000 ? _T_121[63] : _T_121[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_8_io_is_flip = _T_121[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_9_io_in_Re = io_in_9_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_9_io_in_Im = io_in_9_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_9_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_9_io_is_neg = _T_136[62:32] == 31'h3f800000 ? _T_136[63] : _T_136[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_9_io_is_flip = _T_136[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_10_io_in_Re = io_in_10_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_10_io_in_Im = io_in_10_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_10_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_10_io_is_neg = _T_151[62:32] == 31'h3f800000 ? _T_151[63] : _T_151[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_10_io_is_flip = _T_151[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_11_io_in_Re = io_in_11_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_11_io_in_Im = io_in_11_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_11_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_11_io_is_neg = _T_166[62:32] == 31'h3f800000 ? _T_166[63] : _T_166[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_11_io_is_flip = _T_166[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_12_io_in_Re = io_in_12_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_12_io_in_Im = io_in_12_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_12_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_12_io_is_neg = _T_181[62:32] == 31'h3f800000 ? _T_181[63] : _T_181[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_12_io_is_flip = _T_181[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_13_io_in_Re = io_in_13_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_13_io_in_Im = io_in_13_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_13_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_13_io_is_neg = _T_196[62:32] == 31'h3f800000 ? _T_196[63] : _T_196[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_13_io_is_flip = _T_196[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_14_io_in_Re = io_in_14_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_14_io_in_Im = io_in_14_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_14_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_14_io_is_neg = _T_211[62:32] == 31'h3f800000 ? _T_211[63] : _T_211[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_14_io_is_flip = _T_211[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  assign ComplexMULT_SCAL_NOFP_bw32_15_io_in_Re = io_in_15_Re; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_15_io_in_Im = io_in_15_Im; // @[TwidFactorDesigns.scala 86:29]
  assign ComplexMULT_SCAL_NOFP_bw32_15_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 85:32]
  assign ComplexMULT_SCAL_NOFP_bw32_15_io_is_neg = _T_226[62:32] == 31'h3f800000 ? _T_226[63] : _T_226[31]; // @[TwidFactorDesigns.scala 88:125]
  assign ComplexMULT_SCAL_NOFP_bw32_15_io_is_flip = _T_226[62:32] == 31'h3f800000 ? 1'h0 : 1'h1; // @[TwidFactorDesigns.scala 88:125 89:36 96:36]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en) begin // @[TwidFactorDesigns.scala 57:22]
      if (io_in_valid) begin // @[TwidFactorDesigns.scala 58:27]
        value_1 <= _value_T_1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_Re <= ComplexMULT_SCAL_NOFP_bw32_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_Im <= ComplexMULT_SCAL_NOFP_bw32_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_1_Re <= sr_result_regs_r_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_1_Im <= sr_result_regs_r_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_2_Re <= sr_result_regs_r_1_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_2_Im <= sr_result_regs_r_1_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_3_Re <= sr_result_regs_r_2_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_3_Im <= sr_result_regs_r_2_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_4_Re <= sr_result_regs_r_3_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_4_Im <= sr_result_regs_r_3_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_5_Re <= sr_result_regs_r_4_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_5_Im <= sr_result_regs_r_4_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_6_Re <= sr_result_regs_r_5_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_6_Im <= sr_result_regs_r_5_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_7_Re <= sr_result_regs_r_6_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_7_Im <= sr_result_regs_r_6_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_8_Re <= sr_result_regs_r_7_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_8_Im <= sr_result_regs_r_7_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_9_Re <= sr_result_regs_r_8_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_9_Im <= sr_result_regs_r_8_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_10_Re <= sr_result_regs_r_9_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_10_Im <= sr_result_regs_r_9_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_11_Re <= sr_result_regs_r_10_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_11_Im <= sr_result_regs_r_10_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_12_Re <= sr_result_regs_r_11_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_12_Im <= sr_result_regs_r_11_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_13_Re <= sr_result_regs_r_12_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_13_Im <= sr_result_regs_r_12_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_14_Re <= sr_result_regs_r_13_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_14_Im <= sr_result_regs_r_13_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_15_Re <= sr_result_regs_r_14_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_15_Im <= sr_result_regs_r_14_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_16_Re <= sr_result_regs_r_15_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_16_Im <= sr_result_regs_r_15_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_17_Re <= sr_result_regs_r_16_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_17_Im <= sr_result_regs_r_16_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_18_Re <= sr_result_regs_r_17_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_18_Im <= sr_result_regs_r_17_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_19_Re <= sr_result_regs_r_18_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_19_Im <= sr_result_regs_r_18_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_20_Re <= sr_result_regs_r_19_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_20_Im <= sr_result_regs_r_19_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_21_Re <= sr_result_regs_r_20_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_21_Im <= sr_result_regs_r_20_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_22_Re <= sr_result_regs_r_21_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_22_Im <= sr_result_regs_r_21_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_23_Re <= sr_result_regs_r_22_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_23_Im <= sr_result_regs_r_22_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_24_Re <= ComplexMULT_SCAL_NOFP_bw32_1_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_24_Im <= ComplexMULT_SCAL_NOFP_bw32_1_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_25_Re <= sr_result_regs_r_24_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_25_Im <= sr_result_regs_r_24_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_26_Re <= sr_result_regs_r_25_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_26_Im <= sr_result_regs_r_25_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_27_Re <= sr_result_regs_r_26_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_27_Im <= sr_result_regs_r_26_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_28_Re <= sr_result_regs_r_27_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_28_Im <= sr_result_regs_r_27_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_29_Re <= sr_result_regs_r_28_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_29_Im <= sr_result_regs_r_28_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_30_Re <= sr_result_regs_r_29_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_30_Im <= sr_result_regs_r_29_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_31_Re <= sr_result_regs_r_30_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_31_Im <= sr_result_regs_r_30_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_32_Re <= sr_result_regs_r_31_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_32_Im <= sr_result_regs_r_31_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_33_Re <= sr_result_regs_r_32_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_33_Im <= sr_result_regs_r_32_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_34_Re <= sr_result_regs_r_33_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_34_Im <= sr_result_regs_r_33_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_35_Re <= sr_result_regs_r_34_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_35_Im <= sr_result_regs_r_34_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_36_Re <= sr_result_regs_r_35_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_36_Im <= sr_result_regs_r_35_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_37_Re <= sr_result_regs_r_36_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_37_Im <= sr_result_regs_r_36_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_38_Re <= sr_result_regs_r_37_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_38_Im <= sr_result_regs_r_37_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_39_Re <= sr_result_regs_r_38_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_39_Im <= sr_result_regs_r_38_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_40_Re <= sr_result_regs_r_39_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_40_Im <= sr_result_regs_r_39_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_41_Re <= sr_result_regs_r_40_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_41_Im <= sr_result_regs_r_40_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_42_Re <= sr_result_regs_r_41_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_42_Im <= sr_result_regs_r_41_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_43_Re <= sr_result_regs_r_42_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_43_Im <= sr_result_regs_r_42_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_44_Re <= sr_result_regs_r_43_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_44_Im <= sr_result_regs_r_43_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_45_Re <= sr_result_regs_r_44_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_45_Im <= sr_result_regs_r_44_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_46_Re <= sr_result_regs_r_45_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_46_Im <= sr_result_regs_r_45_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_47_Re <= sr_result_regs_r_46_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_47_Im <= sr_result_regs_r_46_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_48_Re <= ComplexMULT_SCAL_NOFP_bw32_2_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_48_Im <= ComplexMULT_SCAL_NOFP_bw32_2_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_49_Re <= sr_result_regs_r_48_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_49_Im <= sr_result_regs_r_48_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_50_Re <= sr_result_regs_r_49_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_50_Im <= sr_result_regs_r_49_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_51_Re <= sr_result_regs_r_50_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_51_Im <= sr_result_regs_r_50_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_52_Re <= sr_result_regs_r_51_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_52_Im <= sr_result_regs_r_51_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_53_Re <= sr_result_regs_r_52_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_53_Im <= sr_result_regs_r_52_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_54_Re <= sr_result_regs_r_53_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_54_Im <= sr_result_regs_r_53_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_55_Re <= sr_result_regs_r_54_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_55_Im <= sr_result_regs_r_54_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_56_Re <= sr_result_regs_r_55_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_56_Im <= sr_result_regs_r_55_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_57_Re <= sr_result_regs_r_56_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_57_Im <= sr_result_regs_r_56_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_58_Re <= sr_result_regs_r_57_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_58_Im <= sr_result_regs_r_57_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_59_Re <= sr_result_regs_r_58_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_59_Im <= sr_result_regs_r_58_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_60_Re <= sr_result_regs_r_59_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_60_Im <= sr_result_regs_r_59_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_61_Re <= sr_result_regs_r_60_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_61_Im <= sr_result_regs_r_60_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_62_Re <= sr_result_regs_r_61_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_62_Im <= sr_result_regs_r_61_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_63_Re <= sr_result_regs_r_62_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_63_Im <= sr_result_regs_r_62_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_64_Re <= sr_result_regs_r_63_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_64_Im <= sr_result_regs_r_63_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_65_Re <= sr_result_regs_r_64_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_65_Im <= sr_result_regs_r_64_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_66_Re <= sr_result_regs_r_65_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_66_Im <= sr_result_regs_r_65_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_67_Re <= sr_result_regs_r_66_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_67_Im <= sr_result_regs_r_66_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_68_Re <= sr_result_regs_r_67_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_68_Im <= sr_result_regs_r_67_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_69_Re <= sr_result_regs_r_68_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_69_Im <= sr_result_regs_r_68_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_70_Re <= sr_result_regs_r_69_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_70_Im <= sr_result_regs_r_69_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_71_Re <= sr_result_regs_r_70_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_71_Im <= sr_result_regs_r_70_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_72_Re <= ComplexMULT_SCAL_NOFP_bw32_3_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_72_Im <= ComplexMULT_SCAL_NOFP_bw32_3_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_73_Re <= sr_result_regs_r_72_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_73_Im <= sr_result_regs_r_72_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_74_Re <= sr_result_regs_r_73_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_74_Im <= sr_result_regs_r_73_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_75_Re <= sr_result_regs_r_74_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_75_Im <= sr_result_regs_r_74_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_76_Re <= sr_result_regs_r_75_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_76_Im <= sr_result_regs_r_75_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_77_Re <= sr_result_regs_r_76_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_77_Im <= sr_result_regs_r_76_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_78_Re <= sr_result_regs_r_77_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_78_Im <= sr_result_regs_r_77_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_79_Re <= sr_result_regs_r_78_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_79_Im <= sr_result_regs_r_78_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_80_Re <= sr_result_regs_r_79_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_80_Im <= sr_result_regs_r_79_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_81_Re <= sr_result_regs_r_80_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_81_Im <= sr_result_regs_r_80_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_82_Re <= sr_result_regs_r_81_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_82_Im <= sr_result_regs_r_81_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_83_Re <= sr_result_regs_r_82_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_83_Im <= sr_result_regs_r_82_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_84_Re <= sr_result_regs_r_83_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_84_Im <= sr_result_regs_r_83_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_85_Re <= sr_result_regs_r_84_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_85_Im <= sr_result_regs_r_84_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_86_Re <= sr_result_regs_r_85_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_86_Im <= sr_result_regs_r_85_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_87_Re <= sr_result_regs_r_86_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_87_Im <= sr_result_regs_r_86_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_88_Re <= sr_result_regs_r_87_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_88_Im <= sr_result_regs_r_87_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_89_Re <= sr_result_regs_r_88_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_89_Im <= sr_result_regs_r_88_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_90_Re <= sr_result_regs_r_89_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_90_Im <= sr_result_regs_r_89_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_91_Re <= sr_result_regs_r_90_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_91_Im <= sr_result_regs_r_90_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_92_Re <= sr_result_regs_r_91_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_92_Im <= sr_result_regs_r_91_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_93_Re <= sr_result_regs_r_92_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_93_Im <= sr_result_regs_r_92_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_94_Re <= sr_result_regs_r_93_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_94_Im <= sr_result_regs_r_93_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_95_Re <= sr_result_regs_r_94_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_95_Im <= sr_result_regs_r_94_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_96_Re <= ComplexMULT_SCAL_NOFP_bw32_4_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_96_Im <= ComplexMULT_SCAL_NOFP_bw32_4_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_97_Re <= sr_result_regs_r_96_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_97_Im <= sr_result_regs_r_96_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_98_Re <= sr_result_regs_r_97_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_98_Im <= sr_result_regs_r_97_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_99_Re <= sr_result_regs_r_98_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_99_Im <= sr_result_regs_r_98_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_100_Re <= sr_result_regs_r_99_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_100_Im <= sr_result_regs_r_99_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_101_Re <= sr_result_regs_r_100_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_101_Im <= sr_result_regs_r_100_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_102_Re <= sr_result_regs_r_101_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_102_Im <= sr_result_regs_r_101_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_103_Re <= sr_result_regs_r_102_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_103_Im <= sr_result_regs_r_102_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_104_Re <= sr_result_regs_r_103_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_104_Im <= sr_result_regs_r_103_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_105_Re <= sr_result_regs_r_104_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_105_Im <= sr_result_regs_r_104_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_106_Re <= sr_result_regs_r_105_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_106_Im <= sr_result_regs_r_105_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_107_Re <= sr_result_regs_r_106_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_107_Im <= sr_result_regs_r_106_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_108_Re <= sr_result_regs_r_107_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_108_Im <= sr_result_regs_r_107_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_109_Re <= sr_result_regs_r_108_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_109_Im <= sr_result_regs_r_108_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_110_Re <= sr_result_regs_r_109_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_110_Im <= sr_result_regs_r_109_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_111_Re <= sr_result_regs_r_110_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_111_Im <= sr_result_regs_r_110_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_112_Re <= sr_result_regs_r_111_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_112_Im <= sr_result_regs_r_111_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_113_Re <= sr_result_regs_r_112_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_113_Im <= sr_result_regs_r_112_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_114_Re <= sr_result_regs_r_113_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_114_Im <= sr_result_regs_r_113_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_115_Re <= sr_result_regs_r_114_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_115_Im <= sr_result_regs_r_114_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_116_Re <= sr_result_regs_r_115_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_116_Im <= sr_result_regs_r_115_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_117_Re <= sr_result_regs_r_116_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_117_Im <= sr_result_regs_r_116_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_118_Re <= sr_result_regs_r_117_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_118_Im <= sr_result_regs_r_117_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_119_Re <= sr_result_regs_r_118_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_119_Im <= sr_result_regs_r_118_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_120_Re <= ComplexMULT_SCAL_NOFP_bw32_5_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_120_Im <= ComplexMULT_SCAL_NOFP_bw32_5_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_121_Re <= sr_result_regs_r_120_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_121_Im <= sr_result_regs_r_120_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_122_Re <= sr_result_regs_r_121_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_122_Im <= sr_result_regs_r_121_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_123_Re <= sr_result_regs_r_122_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_123_Im <= sr_result_regs_r_122_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_124_Re <= sr_result_regs_r_123_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_124_Im <= sr_result_regs_r_123_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_125_Re <= sr_result_regs_r_124_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_125_Im <= sr_result_regs_r_124_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_126_Re <= sr_result_regs_r_125_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_126_Im <= sr_result_regs_r_125_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_127_Re <= sr_result_regs_r_126_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_127_Im <= sr_result_regs_r_126_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_128_Re <= sr_result_regs_r_127_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_128_Im <= sr_result_regs_r_127_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_129_Re <= sr_result_regs_r_128_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_129_Im <= sr_result_regs_r_128_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_130_Re <= sr_result_regs_r_129_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_130_Im <= sr_result_regs_r_129_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_131_Re <= sr_result_regs_r_130_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_131_Im <= sr_result_regs_r_130_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_132_Re <= sr_result_regs_r_131_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_132_Im <= sr_result_regs_r_131_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_133_Re <= sr_result_regs_r_132_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_133_Im <= sr_result_regs_r_132_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_134_Re <= sr_result_regs_r_133_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_134_Im <= sr_result_regs_r_133_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_135_Re <= sr_result_regs_r_134_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_135_Im <= sr_result_regs_r_134_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_136_Re <= sr_result_regs_r_135_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_136_Im <= sr_result_regs_r_135_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_137_Re <= sr_result_regs_r_136_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_137_Im <= sr_result_regs_r_136_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_138_Re <= sr_result_regs_r_137_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_138_Im <= sr_result_regs_r_137_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_139_Re <= sr_result_regs_r_138_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_139_Im <= sr_result_regs_r_138_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_140_Re <= sr_result_regs_r_139_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_140_Im <= sr_result_regs_r_139_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_141_Re <= sr_result_regs_r_140_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_141_Im <= sr_result_regs_r_140_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_142_Re <= sr_result_regs_r_141_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_142_Im <= sr_result_regs_r_141_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_143_Re <= sr_result_regs_r_142_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_143_Im <= sr_result_regs_r_142_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_144_Re <= ComplexMULT_SCAL_NOFP_bw32_6_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_144_Im <= ComplexMULT_SCAL_NOFP_bw32_6_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_145_Re <= sr_result_regs_r_144_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_145_Im <= sr_result_regs_r_144_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_146_Re <= sr_result_regs_r_145_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_146_Im <= sr_result_regs_r_145_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_147_Re <= sr_result_regs_r_146_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_147_Im <= sr_result_regs_r_146_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_148_Re <= sr_result_regs_r_147_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_148_Im <= sr_result_regs_r_147_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_149_Re <= sr_result_regs_r_148_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_149_Im <= sr_result_regs_r_148_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_150_Re <= sr_result_regs_r_149_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_150_Im <= sr_result_regs_r_149_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_151_Re <= sr_result_regs_r_150_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_151_Im <= sr_result_regs_r_150_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_152_Re <= sr_result_regs_r_151_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_152_Im <= sr_result_regs_r_151_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_153_Re <= sr_result_regs_r_152_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_153_Im <= sr_result_regs_r_152_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_154_Re <= sr_result_regs_r_153_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_154_Im <= sr_result_regs_r_153_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_155_Re <= sr_result_regs_r_154_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_155_Im <= sr_result_regs_r_154_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_156_Re <= sr_result_regs_r_155_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_156_Im <= sr_result_regs_r_155_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_157_Re <= sr_result_regs_r_156_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_157_Im <= sr_result_regs_r_156_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_158_Re <= sr_result_regs_r_157_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_158_Im <= sr_result_regs_r_157_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_159_Re <= sr_result_regs_r_158_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_159_Im <= sr_result_regs_r_158_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_160_Re <= sr_result_regs_r_159_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_160_Im <= sr_result_regs_r_159_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_161_Re <= sr_result_regs_r_160_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_161_Im <= sr_result_regs_r_160_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_162_Re <= sr_result_regs_r_161_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_162_Im <= sr_result_regs_r_161_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_163_Re <= sr_result_regs_r_162_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_163_Im <= sr_result_regs_r_162_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_164_Re <= sr_result_regs_r_163_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_164_Im <= sr_result_regs_r_163_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_165_Re <= sr_result_regs_r_164_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_165_Im <= sr_result_regs_r_164_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_166_Re <= sr_result_regs_r_165_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_166_Im <= sr_result_regs_r_165_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_167_Re <= sr_result_regs_r_166_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_167_Im <= sr_result_regs_r_166_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_168_Re <= ComplexMULT_SCAL_NOFP_bw32_7_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_168_Im <= ComplexMULT_SCAL_NOFP_bw32_7_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_169_Re <= sr_result_regs_r_168_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_169_Im <= sr_result_regs_r_168_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_170_Re <= sr_result_regs_r_169_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_170_Im <= sr_result_regs_r_169_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_171_Re <= sr_result_regs_r_170_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_171_Im <= sr_result_regs_r_170_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_172_Re <= sr_result_regs_r_171_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_172_Im <= sr_result_regs_r_171_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_173_Re <= sr_result_regs_r_172_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_173_Im <= sr_result_regs_r_172_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_174_Re <= sr_result_regs_r_173_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_174_Im <= sr_result_regs_r_173_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_175_Re <= sr_result_regs_r_174_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_175_Im <= sr_result_regs_r_174_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_176_Re <= sr_result_regs_r_175_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_176_Im <= sr_result_regs_r_175_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_177_Re <= sr_result_regs_r_176_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_177_Im <= sr_result_regs_r_176_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_178_Re <= sr_result_regs_r_177_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_178_Im <= sr_result_regs_r_177_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_179_Re <= sr_result_regs_r_178_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_179_Im <= sr_result_regs_r_178_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_180_Re <= sr_result_regs_r_179_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_180_Im <= sr_result_regs_r_179_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_181_Re <= sr_result_regs_r_180_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_181_Im <= sr_result_regs_r_180_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_182_Re <= sr_result_regs_r_181_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_182_Im <= sr_result_regs_r_181_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_183_Re <= sr_result_regs_r_182_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_183_Im <= sr_result_regs_r_182_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_184_Re <= sr_result_regs_r_183_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_184_Im <= sr_result_regs_r_183_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_185_Re <= sr_result_regs_r_184_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_185_Im <= sr_result_regs_r_184_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_186_Re <= sr_result_regs_r_185_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_186_Im <= sr_result_regs_r_185_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_187_Re <= sr_result_regs_r_186_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_187_Im <= sr_result_regs_r_186_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_188_Re <= sr_result_regs_r_187_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_188_Im <= sr_result_regs_r_187_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_189_Re <= sr_result_regs_r_188_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_189_Im <= sr_result_regs_r_188_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_190_Re <= sr_result_regs_r_189_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_190_Im <= sr_result_regs_r_189_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_191_Re <= sr_result_regs_r_190_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_191_Im <= sr_result_regs_r_190_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_192_Re <= ComplexMULT_SCAL_NOFP_bw32_8_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_192_Im <= ComplexMULT_SCAL_NOFP_bw32_8_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_193_Re <= sr_result_regs_r_192_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_193_Im <= sr_result_regs_r_192_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_194_Re <= sr_result_regs_r_193_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_194_Im <= sr_result_regs_r_193_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_195_Re <= sr_result_regs_r_194_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_195_Im <= sr_result_regs_r_194_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_196_Re <= sr_result_regs_r_195_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_196_Im <= sr_result_regs_r_195_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_197_Re <= sr_result_regs_r_196_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_197_Im <= sr_result_regs_r_196_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_198_Re <= sr_result_regs_r_197_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_198_Im <= sr_result_regs_r_197_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_199_Re <= sr_result_regs_r_198_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_199_Im <= sr_result_regs_r_198_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_200_Re <= sr_result_regs_r_199_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_200_Im <= sr_result_regs_r_199_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_201_Re <= sr_result_regs_r_200_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_201_Im <= sr_result_regs_r_200_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_202_Re <= sr_result_regs_r_201_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_202_Im <= sr_result_regs_r_201_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_203_Re <= sr_result_regs_r_202_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_203_Im <= sr_result_regs_r_202_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_204_Re <= sr_result_regs_r_203_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_204_Im <= sr_result_regs_r_203_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_205_Re <= sr_result_regs_r_204_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_205_Im <= sr_result_regs_r_204_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_206_Re <= sr_result_regs_r_205_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_206_Im <= sr_result_regs_r_205_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_207_Re <= sr_result_regs_r_206_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_207_Im <= sr_result_regs_r_206_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_208_Re <= sr_result_regs_r_207_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_208_Im <= sr_result_regs_r_207_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_209_Re <= sr_result_regs_r_208_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_209_Im <= sr_result_regs_r_208_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_210_Re <= sr_result_regs_r_209_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_210_Im <= sr_result_regs_r_209_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_211_Re <= sr_result_regs_r_210_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_211_Im <= sr_result_regs_r_210_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_212_Re <= sr_result_regs_r_211_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_212_Im <= sr_result_regs_r_211_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_213_Re <= sr_result_regs_r_212_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_213_Im <= sr_result_regs_r_212_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_214_Re <= sr_result_regs_r_213_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_214_Im <= sr_result_regs_r_213_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_215_Re <= sr_result_regs_r_214_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_215_Im <= sr_result_regs_r_214_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_216_Re <= ComplexMULT_SCAL_NOFP_bw32_9_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_216_Im <= ComplexMULT_SCAL_NOFP_bw32_9_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_217_Re <= sr_result_regs_r_216_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_217_Im <= sr_result_regs_r_216_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_218_Re <= sr_result_regs_r_217_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_218_Im <= sr_result_regs_r_217_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_219_Re <= sr_result_regs_r_218_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_219_Im <= sr_result_regs_r_218_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_220_Re <= sr_result_regs_r_219_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_220_Im <= sr_result_regs_r_219_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_221_Re <= sr_result_regs_r_220_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_221_Im <= sr_result_regs_r_220_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_222_Re <= sr_result_regs_r_221_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_222_Im <= sr_result_regs_r_221_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_223_Re <= sr_result_regs_r_222_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_223_Im <= sr_result_regs_r_222_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_224_Re <= sr_result_regs_r_223_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_224_Im <= sr_result_regs_r_223_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_225_Re <= sr_result_regs_r_224_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_225_Im <= sr_result_regs_r_224_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_226_Re <= sr_result_regs_r_225_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_226_Im <= sr_result_regs_r_225_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_227_Re <= sr_result_regs_r_226_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_227_Im <= sr_result_regs_r_226_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_228_Re <= sr_result_regs_r_227_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_228_Im <= sr_result_regs_r_227_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_229_Re <= sr_result_regs_r_228_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_229_Im <= sr_result_regs_r_228_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_230_Re <= sr_result_regs_r_229_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_230_Im <= sr_result_regs_r_229_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_231_Re <= sr_result_regs_r_230_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_231_Im <= sr_result_regs_r_230_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_232_Re <= sr_result_regs_r_231_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_232_Im <= sr_result_regs_r_231_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_233_Re <= sr_result_regs_r_232_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_233_Im <= sr_result_regs_r_232_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_234_Re <= sr_result_regs_r_233_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_234_Im <= sr_result_regs_r_233_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_235_Re <= sr_result_regs_r_234_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_235_Im <= sr_result_regs_r_234_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_236_Re <= sr_result_regs_r_235_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_236_Im <= sr_result_regs_r_235_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_237_Re <= sr_result_regs_r_236_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_237_Im <= sr_result_regs_r_236_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_238_Re <= sr_result_regs_r_237_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_238_Im <= sr_result_regs_r_237_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_239_Re <= sr_result_regs_r_238_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_239_Im <= sr_result_regs_r_238_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_240_Re <= ComplexMULT_SCAL_NOFP_bw32_10_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_240_Im <= ComplexMULT_SCAL_NOFP_bw32_10_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_241_Re <= sr_result_regs_r_240_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_241_Im <= sr_result_regs_r_240_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_242_Re <= sr_result_regs_r_241_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_242_Im <= sr_result_regs_r_241_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_243_Re <= sr_result_regs_r_242_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_243_Im <= sr_result_regs_r_242_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_244_Re <= sr_result_regs_r_243_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_244_Im <= sr_result_regs_r_243_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_245_Re <= sr_result_regs_r_244_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_245_Im <= sr_result_regs_r_244_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_246_Re <= sr_result_regs_r_245_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_246_Im <= sr_result_regs_r_245_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_247_Re <= sr_result_regs_r_246_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_247_Im <= sr_result_regs_r_246_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_248_Re <= sr_result_regs_r_247_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_248_Im <= sr_result_regs_r_247_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_249_Re <= sr_result_regs_r_248_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_249_Im <= sr_result_regs_r_248_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_250_Re <= sr_result_regs_r_249_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_250_Im <= sr_result_regs_r_249_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_251_Re <= sr_result_regs_r_250_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_251_Im <= sr_result_regs_r_250_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_252_Re <= sr_result_regs_r_251_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_252_Im <= sr_result_regs_r_251_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_253_Re <= sr_result_regs_r_252_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_253_Im <= sr_result_regs_r_252_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_254_Re <= sr_result_regs_r_253_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_254_Im <= sr_result_regs_r_253_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_255_Re <= sr_result_regs_r_254_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_255_Im <= sr_result_regs_r_254_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_256_Re <= sr_result_regs_r_255_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_256_Im <= sr_result_regs_r_255_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_257_Re <= sr_result_regs_r_256_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_257_Im <= sr_result_regs_r_256_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_258_Re <= sr_result_regs_r_257_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_258_Im <= sr_result_regs_r_257_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_259_Re <= sr_result_regs_r_258_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_259_Im <= sr_result_regs_r_258_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_260_Re <= sr_result_regs_r_259_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_260_Im <= sr_result_regs_r_259_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_261_Re <= sr_result_regs_r_260_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_261_Im <= sr_result_regs_r_260_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_262_Re <= sr_result_regs_r_261_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_262_Im <= sr_result_regs_r_261_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_263_Re <= sr_result_regs_r_262_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_263_Im <= sr_result_regs_r_262_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_264_Re <= ComplexMULT_SCAL_NOFP_bw32_11_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_264_Im <= ComplexMULT_SCAL_NOFP_bw32_11_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_265_Re <= sr_result_regs_r_264_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_265_Im <= sr_result_regs_r_264_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_266_Re <= sr_result_regs_r_265_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_266_Im <= sr_result_regs_r_265_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_267_Re <= sr_result_regs_r_266_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_267_Im <= sr_result_regs_r_266_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_268_Re <= sr_result_regs_r_267_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_268_Im <= sr_result_regs_r_267_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_269_Re <= sr_result_regs_r_268_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_269_Im <= sr_result_regs_r_268_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_270_Re <= sr_result_regs_r_269_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_270_Im <= sr_result_regs_r_269_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_271_Re <= sr_result_regs_r_270_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_271_Im <= sr_result_regs_r_270_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_272_Re <= sr_result_regs_r_271_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_272_Im <= sr_result_regs_r_271_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_273_Re <= sr_result_regs_r_272_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_273_Im <= sr_result_regs_r_272_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_274_Re <= sr_result_regs_r_273_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_274_Im <= sr_result_regs_r_273_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_275_Re <= sr_result_regs_r_274_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_275_Im <= sr_result_regs_r_274_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_276_Re <= sr_result_regs_r_275_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_276_Im <= sr_result_regs_r_275_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_277_Re <= sr_result_regs_r_276_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_277_Im <= sr_result_regs_r_276_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_278_Re <= sr_result_regs_r_277_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_278_Im <= sr_result_regs_r_277_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_279_Re <= sr_result_regs_r_278_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_279_Im <= sr_result_regs_r_278_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_280_Re <= sr_result_regs_r_279_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_280_Im <= sr_result_regs_r_279_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_281_Re <= sr_result_regs_r_280_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_281_Im <= sr_result_regs_r_280_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_282_Re <= sr_result_regs_r_281_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_282_Im <= sr_result_regs_r_281_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_283_Re <= sr_result_regs_r_282_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_283_Im <= sr_result_regs_r_282_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_284_Re <= sr_result_regs_r_283_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_284_Im <= sr_result_regs_r_283_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_285_Re <= sr_result_regs_r_284_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_285_Im <= sr_result_regs_r_284_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_286_Re <= sr_result_regs_r_285_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_286_Im <= sr_result_regs_r_285_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_287_Re <= sr_result_regs_r_286_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_287_Im <= sr_result_regs_r_286_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_288_Re <= ComplexMULT_SCAL_NOFP_bw32_12_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_288_Im <= ComplexMULT_SCAL_NOFP_bw32_12_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_289_Re <= sr_result_regs_r_288_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_289_Im <= sr_result_regs_r_288_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_290_Re <= sr_result_regs_r_289_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_290_Im <= sr_result_regs_r_289_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_291_Re <= sr_result_regs_r_290_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_291_Im <= sr_result_regs_r_290_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_292_Re <= sr_result_regs_r_291_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_292_Im <= sr_result_regs_r_291_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_293_Re <= sr_result_regs_r_292_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_293_Im <= sr_result_regs_r_292_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_294_Re <= sr_result_regs_r_293_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_294_Im <= sr_result_regs_r_293_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_295_Re <= sr_result_regs_r_294_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_295_Im <= sr_result_regs_r_294_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_296_Re <= sr_result_regs_r_295_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_296_Im <= sr_result_regs_r_295_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_297_Re <= sr_result_regs_r_296_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_297_Im <= sr_result_regs_r_296_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_298_Re <= sr_result_regs_r_297_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_298_Im <= sr_result_regs_r_297_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_299_Re <= sr_result_regs_r_298_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_299_Im <= sr_result_regs_r_298_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_300_Re <= sr_result_regs_r_299_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_300_Im <= sr_result_regs_r_299_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_301_Re <= sr_result_regs_r_300_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_301_Im <= sr_result_regs_r_300_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_302_Re <= sr_result_regs_r_301_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_302_Im <= sr_result_regs_r_301_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_303_Re <= sr_result_regs_r_302_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_303_Im <= sr_result_regs_r_302_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_304_Re <= sr_result_regs_r_303_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_304_Im <= sr_result_regs_r_303_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_305_Re <= sr_result_regs_r_304_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_305_Im <= sr_result_regs_r_304_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_306_Re <= sr_result_regs_r_305_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_306_Im <= sr_result_regs_r_305_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_307_Re <= sr_result_regs_r_306_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_307_Im <= sr_result_regs_r_306_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_308_Re <= sr_result_regs_r_307_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_308_Im <= sr_result_regs_r_307_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_309_Re <= sr_result_regs_r_308_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_309_Im <= sr_result_regs_r_308_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_310_Re <= sr_result_regs_r_309_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_310_Im <= sr_result_regs_r_309_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_311_Re <= sr_result_regs_r_310_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_311_Im <= sr_result_regs_r_310_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_312_Re <= ComplexMULT_SCAL_NOFP_bw32_13_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_312_Im <= ComplexMULT_SCAL_NOFP_bw32_13_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_313_Re <= sr_result_regs_r_312_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_313_Im <= sr_result_regs_r_312_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_314_Re <= sr_result_regs_r_313_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_314_Im <= sr_result_regs_r_313_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_315_Re <= sr_result_regs_r_314_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_315_Im <= sr_result_regs_r_314_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_316_Re <= sr_result_regs_r_315_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_316_Im <= sr_result_regs_r_315_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_317_Re <= sr_result_regs_r_316_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_317_Im <= sr_result_regs_r_316_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_318_Re <= sr_result_regs_r_317_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_318_Im <= sr_result_regs_r_317_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_319_Re <= sr_result_regs_r_318_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_319_Im <= sr_result_regs_r_318_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_320_Re <= sr_result_regs_r_319_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_320_Im <= sr_result_regs_r_319_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_321_Re <= sr_result_regs_r_320_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_321_Im <= sr_result_regs_r_320_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_322_Re <= sr_result_regs_r_321_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_322_Im <= sr_result_regs_r_321_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_323_Re <= sr_result_regs_r_322_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_323_Im <= sr_result_regs_r_322_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_324_Re <= sr_result_regs_r_323_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_324_Im <= sr_result_regs_r_323_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_325_Re <= sr_result_regs_r_324_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_325_Im <= sr_result_regs_r_324_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_326_Re <= sr_result_regs_r_325_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_326_Im <= sr_result_regs_r_325_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_327_Re <= sr_result_regs_r_326_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_327_Im <= sr_result_regs_r_326_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_328_Re <= sr_result_regs_r_327_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_328_Im <= sr_result_regs_r_327_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_329_Re <= sr_result_regs_r_328_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_329_Im <= sr_result_regs_r_328_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_330_Re <= sr_result_regs_r_329_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_330_Im <= sr_result_regs_r_329_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_331_Re <= sr_result_regs_r_330_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_331_Im <= sr_result_regs_r_330_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_332_Re <= sr_result_regs_r_331_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_332_Im <= sr_result_regs_r_331_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_333_Re <= sr_result_regs_r_332_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_333_Im <= sr_result_regs_r_332_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_334_Re <= sr_result_regs_r_333_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_334_Im <= sr_result_regs_r_333_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_335_Re <= sr_result_regs_r_334_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_335_Im <= sr_result_regs_r_334_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_336_Re <= ComplexMULT_SCAL_NOFP_bw32_14_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_336_Im <= ComplexMULT_SCAL_NOFP_bw32_14_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_337_Re <= sr_result_regs_r_336_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_337_Im <= sr_result_regs_r_336_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_338_Re <= sr_result_regs_r_337_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_338_Im <= sr_result_regs_r_337_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_339_Re <= sr_result_regs_r_338_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_339_Im <= sr_result_regs_r_338_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_340_Re <= sr_result_regs_r_339_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_340_Im <= sr_result_regs_r_339_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_341_Re <= sr_result_regs_r_340_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_341_Im <= sr_result_regs_r_340_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_342_Re <= sr_result_regs_r_341_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_342_Im <= sr_result_regs_r_341_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_343_Re <= sr_result_regs_r_342_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_343_Im <= sr_result_regs_r_342_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_344_Re <= sr_result_regs_r_343_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_344_Im <= sr_result_regs_r_343_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_345_Re <= sr_result_regs_r_344_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_345_Im <= sr_result_regs_r_344_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_346_Re <= sr_result_regs_r_345_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_346_Im <= sr_result_regs_r_345_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_347_Re <= sr_result_regs_r_346_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_347_Im <= sr_result_regs_r_346_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_348_Re <= sr_result_regs_r_347_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_348_Im <= sr_result_regs_r_347_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_349_Re <= sr_result_regs_r_348_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_349_Im <= sr_result_regs_r_348_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_350_Re <= sr_result_regs_r_349_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_350_Im <= sr_result_regs_r_349_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_351_Re <= sr_result_regs_r_350_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_351_Im <= sr_result_regs_r_350_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_352_Re <= sr_result_regs_r_351_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_352_Im <= sr_result_regs_r_351_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_353_Re <= sr_result_regs_r_352_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_353_Im <= sr_result_regs_r_352_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_354_Re <= sr_result_regs_r_353_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_354_Im <= sr_result_regs_r_353_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_355_Re <= sr_result_regs_r_354_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_355_Im <= sr_result_regs_r_354_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_356_Re <= sr_result_regs_r_355_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_356_Im <= sr_result_regs_r_355_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_357_Re <= sr_result_regs_r_356_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_357_Im <= sr_result_regs_r_356_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_358_Re <= sr_result_regs_r_357_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_358_Im <= sr_result_regs_r_357_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_359_Re <= sr_result_regs_r_358_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_359_Im <= sr_result_regs_r_358_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_360_Re <= ComplexMULT_SCAL_NOFP_bw32_15_io_out_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_360_Im <= ComplexMULT_SCAL_NOFP_bw32_15_io_out_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_361_Re <= sr_result_regs_r_360_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_361_Im <= sr_result_regs_r_360_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_362_Re <= sr_result_regs_r_361_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_362_Im <= sr_result_regs_r_361_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_363_Re <= sr_result_regs_r_362_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_363_Im <= sr_result_regs_r_362_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_364_Re <= sr_result_regs_r_363_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_364_Im <= sr_result_regs_r_363_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_365_Re <= sr_result_regs_r_364_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_365_Im <= sr_result_regs_r_364_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_366_Re <= sr_result_regs_r_365_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_366_Im <= sr_result_regs_r_365_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_367_Re <= sr_result_regs_r_366_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_367_Im <= sr_result_regs_r_366_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_368_Re <= sr_result_regs_r_367_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_368_Im <= sr_result_regs_r_367_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_369_Re <= sr_result_regs_r_368_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_369_Im <= sr_result_regs_r_368_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_370_Re <= sr_result_regs_r_369_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_370_Im <= sr_result_regs_r_369_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_371_Re <= sr_result_regs_r_370_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_371_Im <= sr_result_regs_r_370_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_372_Re <= sr_result_regs_r_371_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_372_Im <= sr_result_regs_r_371_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_373_Re <= sr_result_regs_r_372_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_373_Im <= sr_result_regs_r_372_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_374_Re <= sr_result_regs_r_373_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_374_Im <= sr_result_regs_r_373_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_375_Re <= sr_result_regs_r_374_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_375_Im <= sr_result_regs_r_374_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_376_Re <= sr_result_regs_r_375_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_376_Im <= sr_result_regs_r_375_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_377_Re <= sr_result_regs_r_376_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_377_Im <= sr_result_regs_r_376_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_378_Re <= sr_result_regs_r_377_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_378_Im <= sr_result_regs_r_377_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_379_Re <= sr_result_regs_r_378_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_379_Im <= sr_result_regs_r_378_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_380_Re <= sr_result_regs_r_379_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_380_Im <= sr_result_regs_r_379_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_381_Re <= sr_result_regs_r_380_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_381_Im <= sr_result_regs_r_380_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_382_Re <= sr_result_regs_r_381_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_382_Im <= sr_result_regs_r_381_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_383_Re <= sr_result_regs_r_382_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      sr_result_regs_r_383_Im <= sr_result_regs_r_382_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r <= io_in_valid; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_1 <= io_out_valid_r; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_2 <= io_out_valid_r_1; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_3 <= io_out_valid_r_2; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_4 <= io_out_valid_r_3; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_5 <= io_out_valid_r_4; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_6 <= io_out_valid_r_5; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_7 <= io_out_valid_r_6; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_8 <= io_out_valid_r_7; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_9 <= io_out_valid_r_8; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_10 <= io_out_valid_r_9; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_11 <= io_out_valid_r_10; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_12 <= io_out_valid_r_11; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_13 <= io_out_valid_r_12; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_14 <= io_out_valid_r_13; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_15 <= io_out_valid_r_14; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_16 <= io_out_valid_r_15; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_17 <= io_out_valid_r_16; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_18 <= io_out_valid_r_17; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_19 <= io_out_valid_r_18; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_20 <= io_out_valid_r_19; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_21 <= io_out_valid_r_20; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_22 <= io_out_valid_r_21; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_23 <= io_out_valid_r_22; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sr_result_regs_r_Re = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  sr_result_regs_r_Im = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  sr_result_regs_r_1_Re = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  sr_result_regs_r_1_Im = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  sr_result_regs_r_2_Re = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  sr_result_regs_r_2_Im = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  sr_result_regs_r_3_Re = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  sr_result_regs_r_3_Im = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  sr_result_regs_r_4_Re = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  sr_result_regs_r_4_Im = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  sr_result_regs_r_5_Re = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  sr_result_regs_r_5_Im = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  sr_result_regs_r_6_Re = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  sr_result_regs_r_6_Im = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  sr_result_regs_r_7_Re = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  sr_result_regs_r_7_Im = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  sr_result_regs_r_8_Re = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  sr_result_regs_r_8_Im = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  sr_result_regs_r_9_Re = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  sr_result_regs_r_9_Im = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  sr_result_regs_r_10_Re = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  sr_result_regs_r_10_Im = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  sr_result_regs_r_11_Re = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  sr_result_regs_r_11_Im = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  sr_result_regs_r_12_Re = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  sr_result_regs_r_12_Im = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  sr_result_regs_r_13_Re = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  sr_result_regs_r_13_Im = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  sr_result_regs_r_14_Re = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  sr_result_regs_r_14_Im = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  sr_result_regs_r_15_Re = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  sr_result_regs_r_15_Im = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  sr_result_regs_r_16_Re = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  sr_result_regs_r_16_Im = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  sr_result_regs_r_17_Re = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  sr_result_regs_r_17_Im = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  sr_result_regs_r_18_Re = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  sr_result_regs_r_18_Im = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  sr_result_regs_r_19_Re = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  sr_result_regs_r_19_Im = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  sr_result_regs_r_20_Re = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  sr_result_regs_r_20_Im = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  sr_result_regs_r_21_Re = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  sr_result_regs_r_21_Im = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  sr_result_regs_r_22_Re = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  sr_result_regs_r_22_Im = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  sr_result_regs_r_23_Re = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  sr_result_regs_r_23_Im = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  sr_result_regs_r_24_Re = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  sr_result_regs_r_24_Im = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  sr_result_regs_r_25_Re = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  sr_result_regs_r_25_Im = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  sr_result_regs_r_26_Re = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  sr_result_regs_r_26_Im = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  sr_result_regs_r_27_Re = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  sr_result_regs_r_27_Im = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  sr_result_regs_r_28_Re = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  sr_result_regs_r_28_Im = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  sr_result_regs_r_29_Re = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  sr_result_regs_r_29_Im = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  sr_result_regs_r_30_Re = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  sr_result_regs_r_30_Im = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  sr_result_regs_r_31_Re = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  sr_result_regs_r_31_Im = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  sr_result_regs_r_32_Re = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  sr_result_regs_r_32_Im = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sr_result_regs_r_33_Re = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  sr_result_regs_r_33_Im = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  sr_result_regs_r_34_Re = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  sr_result_regs_r_34_Im = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  sr_result_regs_r_35_Re = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  sr_result_regs_r_35_Im = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  sr_result_regs_r_36_Re = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  sr_result_regs_r_36_Im = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  sr_result_regs_r_37_Re = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  sr_result_regs_r_37_Im = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  sr_result_regs_r_38_Re = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  sr_result_regs_r_38_Im = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  sr_result_regs_r_39_Re = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  sr_result_regs_r_39_Im = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  sr_result_regs_r_40_Re = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  sr_result_regs_r_40_Im = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  sr_result_regs_r_41_Re = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  sr_result_regs_r_41_Im = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  sr_result_regs_r_42_Re = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  sr_result_regs_r_42_Im = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  sr_result_regs_r_43_Re = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  sr_result_regs_r_43_Im = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  sr_result_regs_r_44_Re = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  sr_result_regs_r_44_Im = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  sr_result_regs_r_45_Re = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  sr_result_regs_r_45_Im = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  sr_result_regs_r_46_Re = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  sr_result_regs_r_46_Im = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  sr_result_regs_r_47_Re = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  sr_result_regs_r_47_Im = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  sr_result_regs_r_48_Re = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  sr_result_regs_r_48_Im = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  sr_result_regs_r_49_Re = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  sr_result_regs_r_49_Im = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  sr_result_regs_r_50_Re = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  sr_result_regs_r_50_Im = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  sr_result_regs_r_51_Re = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  sr_result_regs_r_51_Im = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  sr_result_regs_r_52_Re = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  sr_result_regs_r_52_Im = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  sr_result_regs_r_53_Re = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  sr_result_regs_r_53_Im = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  sr_result_regs_r_54_Re = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  sr_result_regs_r_54_Im = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  sr_result_regs_r_55_Re = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  sr_result_regs_r_55_Im = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  sr_result_regs_r_56_Re = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  sr_result_regs_r_56_Im = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  sr_result_regs_r_57_Re = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  sr_result_regs_r_57_Im = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  sr_result_regs_r_58_Re = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  sr_result_regs_r_58_Im = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  sr_result_regs_r_59_Re = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  sr_result_regs_r_59_Im = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  sr_result_regs_r_60_Re = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  sr_result_regs_r_60_Im = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  sr_result_regs_r_61_Re = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  sr_result_regs_r_61_Im = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  sr_result_regs_r_62_Re = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  sr_result_regs_r_62_Im = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  sr_result_regs_r_63_Re = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  sr_result_regs_r_63_Im = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  sr_result_regs_r_64_Re = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  sr_result_regs_r_64_Im = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  sr_result_regs_r_65_Re = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  sr_result_regs_r_65_Im = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  sr_result_regs_r_66_Re = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  sr_result_regs_r_66_Im = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  sr_result_regs_r_67_Re = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  sr_result_regs_r_67_Im = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  sr_result_regs_r_68_Re = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  sr_result_regs_r_68_Im = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  sr_result_regs_r_69_Re = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  sr_result_regs_r_69_Im = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  sr_result_regs_r_70_Re = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  sr_result_regs_r_70_Im = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  sr_result_regs_r_71_Re = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  sr_result_regs_r_71_Im = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  sr_result_regs_r_72_Re = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  sr_result_regs_r_72_Im = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  sr_result_regs_r_73_Re = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  sr_result_regs_r_73_Im = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  sr_result_regs_r_74_Re = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  sr_result_regs_r_74_Im = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  sr_result_regs_r_75_Re = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  sr_result_regs_r_75_Im = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  sr_result_regs_r_76_Re = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  sr_result_regs_r_76_Im = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  sr_result_regs_r_77_Re = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  sr_result_regs_r_77_Im = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  sr_result_regs_r_78_Re = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  sr_result_regs_r_78_Im = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  sr_result_regs_r_79_Re = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  sr_result_regs_r_79_Im = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  sr_result_regs_r_80_Re = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  sr_result_regs_r_80_Im = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  sr_result_regs_r_81_Re = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  sr_result_regs_r_81_Im = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  sr_result_regs_r_82_Re = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  sr_result_regs_r_82_Im = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  sr_result_regs_r_83_Re = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  sr_result_regs_r_83_Im = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  sr_result_regs_r_84_Re = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  sr_result_regs_r_84_Im = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  sr_result_regs_r_85_Re = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  sr_result_regs_r_85_Im = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  sr_result_regs_r_86_Re = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  sr_result_regs_r_86_Im = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  sr_result_regs_r_87_Re = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  sr_result_regs_r_87_Im = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  sr_result_regs_r_88_Re = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  sr_result_regs_r_88_Im = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  sr_result_regs_r_89_Re = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  sr_result_regs_r_89_Im = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  sr_result_regs_r_90_Re = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  sr_result_regs_r_90_Im = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  sr_result_regs_r_91_Re = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  sr_result_regs_r_91_Im = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  sr_result_regs_r_92_Re = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  sr_result_regs_r_92_Im = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  sr_result_regs_r_93_Re = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  sr_result_regs_r_93_Im = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  sr_result_regs_r_94_Re = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  sr_result_regs_r_94_Im = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  sr_result_regs_r_95_Re = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  sr_result_regs_r_95_Im = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  sr_result_regs_r_96_Re = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  sr_result_regs_r_96_Im = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  sr_result_regs_r_97_Re = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  sr_result_regs_r_97_Im = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  sr_result_regs_r_98_Re = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  sr_result_regs_r_98_Im = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  sr_result_regs_r_99_Re = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  sr_result_regs_r_99_Im = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  sr_result_regs_r_100_Re = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  sr_result_regs_r_100_Im = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  sr_result_regs_r_101_Re = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  sr_result_regs_r_101_Im = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  sr_result_regs_r_102_Re = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  sr_result_regs_r_102_Im = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  sr_result_regs_r_103_Re = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  sr_result_regs_r_103_Im = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  sr_result_regs_r_104_Re = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  sr_result_regs_r_104_Im = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  sr_result_regs_r_105_Re = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  sr_result_regs_r_105_Im = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  sr_result_regs_r_106_Re = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  sr_result_regs_r_106_Im = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  sr_result_regs_r_107_Re = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  sr_result_regs_r_107_Im = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  sr_result_regs_r_108_Re = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  sr_result_regs_r_108_Im = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  sr_result_regs_r_109_Re = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  sr_result_regs_r_109_Im = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  sr_result_regs_r_110_Re = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  sr_result_regs_r_110_Im = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  sr_result_regs_r_111_Re = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  sr_result_regs_r_111_Im = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  sr_result_regs_r_112_Re = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  sr_result_regs_r_112_Im = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  sr_result_regs_r_113_Re = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  sr_result_regs_r_113_Im = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  sr_result_regs_r_114_Re = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  sr_result_regs_r_114_Im = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  sr_result_regs_r_115_Re = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  sr_result_regs_r_115_Im = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  sr_result_regs_r_116_Re = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  sr_result_regs_r_116_Im = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  sr_result_regs_r_117_Re = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  sr_result_regs_r_117_Im = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  sr_result_regs_r_118_Re = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  sr_result_regs_r_118_Im = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  sr_result_regs_r_119_Re = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  sr_result_regs_r_119_Im = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  sr_result_regs_r_120_Re = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  sr_result_regs_r_120_Im = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  sr_result_regs_r_121_Re = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  sr_result_regs_r_121_Im = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  sr_result_regs_r_122_Re = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  sr_result_regs_r_122_Im = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  sr_result_regs_r_123_Re = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  sr_result_regs_r_123_Im = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  sr_result_regs_r_124_Re = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  sr_result_regs_r_124_Im = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  sr_result_regs_r_125_Re = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  sr_result_regs_r_125_Im = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  sr_result_regs_r_126_Re = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  sr_result_regs_r_126_Im = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  sr_result_regs_r_127_Re = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  sr_result_regs_r_127_Im = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  sr_result_regs_r_128_Re = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  sr_result_regs_r_128_Im = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  sr_result_regs_r_129_Re = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  sr_result_regs_r_129_Im = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  sr_result_regs_r_130_Re = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  sr_result_regs_r_130_Im = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  sr_result_regs_r_131_Re = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  sr_result_regs_r_131_Im = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  sr_result_regs_r_132_Re = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  sr_result_regs_r_132_Im = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  sr_result_regs_r_133_Re = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  sr_result_regs_r_133_Im = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  sr_result_regs_r_134_Re = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  sr_result_regs_r_134_Im = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  sr_result_regs_r_135_Re = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  sr_result_regs_r_135_Im = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  sr_result_regs_r_136_Re = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  sr_result_regs_r_136_Im = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  sr_result_regs_r_137_Re = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  sr_result_regs_r_137_Im = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  sr_result_regs_r_138_Re = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  sr_result_regs_r_138_Im = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  sr_result_regs_r_139_Re = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  sr_result_regs_r_139_Im = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  sr_result_regs_r_140_Re = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  sr_result_regs_r_140_Im = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  sr_result_regs_r_141_Re = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  sr_result_regs_r_141_Im = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  sr_result_regs_r_142_Re = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  sr_result_regs_r_142_Im = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  sr_result_regs_r_143_Re = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  sr_result_regs_r_143_Im = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  sr_result_regs_r_144_Re = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  sr_result_regs_r_144_Im = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  sr_result_regs_r_145_Re = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  sr_result_regs_r_145_Im = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  sr_result_regs_r_146_Re = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  sr_result_regs_r_146_Im = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  sr_result_regs_r_147_Re = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  sr_result_regs_r_147_Im = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  sr_result_regs_r_148_Re = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  sr_result_regs_r_148_Im = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  sr_result_regs_r_149_Re = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  sr_result_regs_r_149_Im = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  sr_result_regs_r_150_Re = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  sr_result_regs_r_150_Im = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  sr_result_regs_r_151_Re = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  sr_result_regs_r_151_Im = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  sr_result_regs_r_152_Re = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  sr_result_regs_r_152_Im = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  sr_result_regs_r_153_Re = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  sr_result_regs_r_153_Im = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  sr_result_regs_r_154_Re = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  sr_result_regs_r_154_Im = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  sr_result_regs_r_155_Re = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  sr_result_regs_r_155_Im = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  sr_result_regs_r_156_Re = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  sr_result_regs_r_156_Im = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  sr_result_regs_r_157_Re = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  sr_result_regs_r_157_Im = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  sr_result_regs_r_158_Re = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  sr_result_regs_r_158_Im = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  sr_result_regs_r_159_Re = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  sr_result_regs_r_159_Im = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  sr_result_regs_r_160_Re = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  sr_result_regs_r_160_Im = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  sr_result_regs_r_161_Re = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  sr_result_regs_r_161_Im = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  sr_result_regs_r_162_Re = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  sr_result_regs_r_162_Im = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  sr_result_regs_r_163_Re = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  sr_result_regs_r_163_Im = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  sr_result_regs_r_164_Re = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  sr_result_regs_r_164_Im = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  sr_result_regs_r_165_Re = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  sr_result_regs_r_165_Im = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  sr_result_regs_r_166_Re = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  sr_result_regs_r_166_Im = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  sr_result_regs_r_167_Re = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  sr_result_regs_r_167_Im = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  sr_result_regs_r_168_Re = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  sr_result_regs_r_168_Im = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  sr_result_regs_r_169_Re = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  sr_result_regs_r_169_Im = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  sr_result_regs_r_170_Re = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  sr_result_regs_r_170_Im = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  sr_result_regs_r_171_Re = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  sr_result_regs_r_171_Im = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  sr_result_regs_r_172_Re = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  sr_result_regs_r_172_Im = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  sr_result_regs_r_173_Re = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  sr_result_regs_r_173_Im = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  sr_result_regs_r_174_Re = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  sr_result_regs_r_174_Im = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  sr_result_regs_r_175_Re = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  sr_result_regs_r_175_Im = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  sr_result_regs_r_176_Re = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  sr_result_regs_r_176_Im = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  sr_result_regs_r_177_Re = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  sr_result_regs_r_177_Im = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  sr_result_regs_r_178_Re = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  sr_result_regs_r_178_Im = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  sr_result_regs_r_179_Re = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  sr_result_regs_r_179_Im = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  sr_result_regs_r_180_Re = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  sr_result_regs_r_180_Im = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  sr_result_regs_r_181_Re = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  sr_result_regs_r_181_Im = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  sr_result_regs_r_182_Re = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  sr_result_regs_r_182_Im = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  sr_result_regs_r_183_Re = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  sr_result_regs_r_183_Im = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  sr_result_regs_r_184_Re = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  sr_result_regs_r_184_Im = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  sr_result_regs_r_185_Re = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  sr_result_regs_r_185_Im = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  sr_result_regs_r_186_Re = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  sr_result_regs_r_186_Im = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  sr_result_regs_r_187_Re = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  sr_result_regs_r_187_Im = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  sr_result_regs_r_188_Re = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  sr_result_regs_r_188_Im = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  sr_result_regs_r_189_Re = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  sr_result_regs_r_189_Im = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  sr_result_regs_r_190_Re = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  sr_result_regs_r_190_Im = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  sr_result_regs_r_191_Re = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  sr_result_regs_r_191_Im = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  sr_result_regs_r_192_Re = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  sr_result_regs_r_192_Im = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  sr_result_regs_r_193_Re = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  sr_result_regs_r_193_Im = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  sr_result_regs_r_194_Re = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  sr_result_regs_r_194_Im = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  sr_result_regs_r_195_Re = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  sr_result_regs_r_195_Im = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  sr_result_regs_r_196_Re = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  sr_result_regs_r_196_Im = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  sr_result_regs_r_197_Re = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  sr_result_regs_r_197_Im = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  sr_result_regs_r_198_Re = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  sr_result_regs_r_198_Im = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  sr_result_regs_r_199_Re = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  sr_result_regs_r_199_Im = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  sr_result_regs_r_200_Re = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  sr_result_regs_r_200_Im = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  sr_result_regs_r_201_Re = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  sr_result_regs_r_201_Im = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  sr_result_regs_r_202_Re = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  sr_result_regs_r_202_Im = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  sr_result_regs_r_203_Re = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  sr_result_regs_r_203_Im = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  sr_result_regs_r_204_Re = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  sr_result_regs_r_204_Im = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  sr_result_regs_r_205_Re = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  sr_result_regs_r_205_Im = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  sr_result_regs_r_206_Re = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  sr_result_regs_r_206_Im = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  sr_result_regs_r_207_Re = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  sr_result_regs_r_207_Im = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  sr_result_regs_r_208_Re = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  sr_result_regs_r_208_Im = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  sr_result_regs_r_209_Re = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  sr_result_regs_r_209_Im = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  sr_result_regs_r_210_Re = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  sr_result_regs_r_210_Im = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  sr_result_regs_r_211_Re = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  sr_result_regs_r_211_Im = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  sr_result_regs_r_212_Re = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  sr_result_regs_r_212_Im = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  sr_result_regs_r_213_Re = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  sr_result_regs_r_213_Im = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  sr_result_regs_r_214_Re = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  sr_result_regs_r_214_Im = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  sr_result_regs_r_215_Re = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  sr_result_regs_r_215_Im = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  sr_result_regs_r_216_Re = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  sr_result_regs_r_216_Im = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  sr_result_regs_r_217_Re = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  sr_result_regs_r_217_Im = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  sr_result_regs_r_218_Re = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  sr_result_regs_r_218_Im = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  sr_result_regs_r_219_Re = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  sr_result_regs_r_219_Im = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  sr_result_regs_r_220_Re = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  sr_result_regs_r_220_Im = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  sr_result_regs_r_221_Re = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  sr_result_regs_r_221_Im = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  sr_result_regs_r_222_Re = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  sr_result_regs_r_222_Im = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  sr_result_regs_r_223_Re = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  sr_result_regs_r_223_Im = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  sr_result_regs_r_224_Re = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  sr_result_regs_r_224_Im = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  sr_result_regs_r_225_Re = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  sr_result_regs_r_225_Im = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  sr_result_regs_r_226_Re = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  sr_result_regs_r_226_Im = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  sr_result_regs_r_227_Re = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  sr_result_regs_r_227_Im = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  sr_result_regs_r_228_Re = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  sr_result_regs_r_228_Im = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  sr_result_regs_r_229_Re = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  sr_result_regs_r_229_Im = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  sr_result_regs_r_230_Re = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  sr_result_regs_r_230_Im = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  sr_result_regs_r_231_Re = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  sr_result_regs_r_231_Im = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  sr_result_regs_r_232_Re = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  sr_result_regs_r_232_Im = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  sr_result_regs_r_233_Re = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  sr_result_regs_r_233_Im = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  sr_result_regs_r_234_Re = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  sr_result_regs_r_234_Im = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  sr_result_regs_r_235_Re = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  sr_result_regs_r_235_Im = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  sr_result_regs_r_236_Re = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  sr_result_regs_r_236_Im = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  sr_result_regs_r_237_Re = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  sr_result_regs_r_237_Im = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  sr_result_regs_r_238_Re = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  sr_result_regs_r_238_Im = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  sr_result_regs_r_239_Re = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  sr_result_regs_r_239_Im = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  sr_result_regs_r_240_Re = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  sr_result_regs_r_240_Im = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  sr_result_regs_r_241_Re = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  sr_result_regs_r_241_Im = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  sr_result_regs_r_242_Re = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  sr_result_regs_r_242_Im = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  sr_result_regs_r_243_Re = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  sr_result_regs_r_243_Im = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  sr_result_regs_r_244_Re = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  sr_result_regs_r_244_Im = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  sr_result_regs_r_245_Re = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  sr_result_regs_r_245_Im = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  sr_result_regs_r_246_Re = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  sr_result_regs_r_246_Im = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  sr_result_regs_r_247_Re = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  sr_result_regs_r_247_Im = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  sr_result_regs_r_248_Re = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  sr_result_regs_r_248_Im = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  sr_result_regs_r_249_Re = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  sr_result_regs_r_249_Im = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  sr_result_regs_r_250_Re = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  sr_result_regs_r_250_Im = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  sr_result_regs_r_251_Re = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  sr_result_regs_r_251_Im = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  sr_result_regs_r_252_Re = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  sr_result_regs_r_252_Im = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  sr_result_regs_r_253_Re = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  sr_result_regs_r_253_Im = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  sr_result_regs_r_254_Re = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  sr_result_regs_r_254_Im = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  sr_result_regs_r_255_Re = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  sr_result_regs_r_255_Im = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  sr_result_regs_r_256_Re = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  sr_result_regs_r_256_Im = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  sr_result_regs_r_257_Re = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  sr_result_regs_r_257_Im = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  sr_result_regs_r_258_Re = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  sr_result_regs_r_258_Im = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  sr_result_regs_r_259_Re = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  sr_result_regs_r_259_Im = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  sr_result_regs_r_260_Re = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  sr_result_regs_r_260_Im = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  sr_result_regs_r_261_Re = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  sr_result_regs_r_261_Im = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  sr_result_regs_r_262_Re = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  sr_result_regs_r_262_Im = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  sr_result_regs_r_263_Re = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  sr_result_regs_r_263_Im = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  sr_result_regs_r_264_Re = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  sr_result_regs_r_264_Im = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  sr_result_regs_r_265_Re = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  sr_result_regs_r_265_Im = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  sr_result_regs_r_266_Re = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  sr_result_regs_r_266_Im = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  sr_result_regs_r_267_Re = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  sr_result_regs_r_267_Im = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  sr_result_regs_r_268_Re = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  sr_result_regs_r_268_Im = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  sr_result_regs_r_269_Re = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  sr_result_regs_r_269_Im = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  sr_result_regs_r_270_Re = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  sr_result_regs_r_270_Im = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  sr_result_regs_r_271_Re = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  sr_result_regs_r_271_Im = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  sr_result_regs_r_272_Re = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  sr_result_regs_r_272_Im = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  sr_result_regs_r_273_Re = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  sr_result_regs_r_273_Im = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  sr_result_regs_r_274_Re = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  sr_result_regs_r_274_Im = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  sr_result_regs_r_275_Re = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  sr_result_regs_r_275_Im = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  sr_result_regs_r_276_Re = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  sr_result_regs_r_276_Im = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  sr_result_regs_r_277_Re = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  sr_result_regs_r_277_Im = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  sr_result_regs_r_278_Re = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  sr_result_regs_r_278_Im = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  sr_result_regs_r_279_Re = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  sr_result_regs_r_279_Im = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  sr_result_regs_r_280_Re = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  sr_result_regs_r_280_Im = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  sr_result_regs_r_281_Re = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  sr_result_regs_r_281_Im = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  sr_result_regs_r_282_Re = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  sr_result_regs_r_282_Im = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  sr_result_regs_r_283_Re = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  sr_result_regs_r_283_Im = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  sr_result_regs_r_284_Re = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  sr_result_regs_r_284_Im = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  sr_result_regs_r_285_Re = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  sr_result_regs_r_285_Im = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  sr_result_regs_r_286_Re = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  sr_result_regs_r_286_Im = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  sr_result_regs_r_287_Re = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  sr_result_regs_r_287_Im = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  sr_result_regs_r_288_Re = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  sr_result_regs_r_288_Im = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  sr_result_regs_r_289_Re = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  sr_result_regs_r_289_Im = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  sr_result_regs_r_290_Re = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  sr_result_regs_r_290_Im = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  sr_result_regs_r_291_Re = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  sr_result_regs_r_291_Im = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  sr_result_regs_r_292_Re = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  sr_result_regs_r_292_Im = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  sr_result_regs_r_293_Re = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  sr_result_regs_r_293_Im = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  sr_result_regs_r_294_Re = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  sr_result_regs_r_294_Im = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  sr_result_regs_r_295_Re = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  sr_result_regs_r_295_Im = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  sr_result_regs_r_296_Re = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  sr_result_regs_r_296_Im = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  sr_result_regs_r_297_Re = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  sr_result_regs_r_297_Im = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  sr_result_regs_r_298_Re = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  sr_result_regs_r_298_Im = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  sr_result_regs_r_299_Re = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  sr_result_regs_r_299_Im = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  sr_result_regs_r_300_Re = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  sr_result_regs_r_300_Im = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  sr_result_regs_r_301_Re = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  sr_result_regs_r_301_Im = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  sr_result_regs_r_302_Re = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  sr_result_regs_r_302_Im = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  sr_result_regs_r_303_Re = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  sr_result_regs_r_303_Im = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  sr_result_regs_r_304_Re = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  sr_result_regs_r_304_Im = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  sr_result_regs_r_305_Re = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  sr_result_regs_r_305_Im = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  sr_result_regs_r_306_Re = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  sr_result_regs_r_306_Im = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  sr_result_regs_r_307_Re = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  sr_result_regs_r_307_Im = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  sr_result_regs_r_308_Re = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  sr_result_regs_r_308_Im = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  sr_result_regs_r_309_Re = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  sr_result_regs_r_309_Im = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  sr_result_regs_r_310_Re = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  sr_result_regs_r_310_Im = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  sr_result_regs_r_311_Re = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  sr_result_regs_r_311_Im = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  sr_result_regs_r_312_Re = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  sr_result_regs_r_312_Im = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  sr_result_regs_r_313_Re = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  sr_result_regs_r_313_Im = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  sr_result_regs_r_314_Re = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  sr_result_regs_r_314_Im = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  sr_result_regs_r_315_Re = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  sr_result_regs_r_315_Im = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  sr_result_regs_r_316_Re = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  sr_result_regs_r_316_Im = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  sr_result_regs_r_317_Re = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  sr_result_regs_r_317_Im = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  sr_result_regs_r_318_Re = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  sr_result_regs_r_318_Im = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  sr_result_regs_r_319_Re = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  sr_result_regs_r_319_Im = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  sr_result_regs_r_320_Re = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  sr_result_regs_r_320_Im = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  sr_result_regs_r_321_Re = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  sr_result_regs_r_321_Im = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  sr_result_regs_r_322_Re = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  sr_result_regs_r_322_Im = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  sr_result_regs_r_323_Re = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  sr_result_regs_r_323_Im = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  sr_result_regs_r_324_Re = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  sr_result_regs_r_324_Im = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  sr_result_regs_r_325_Re = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  sr_result_regs_r_325_Im = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  sr_result_regs_r_326_Re = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  sr_result_regs_r_326_Im = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  sr_result_regs_r_327_Re = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  sr_result_regs_r_327_Im = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  sr_result_regs_r_328_Re = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  sr_result_regs_r_328_Im = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  sr_result_regs_r_329_Re = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  sr_result_regs_r_329_Im = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  sr_result_regs_r_330_Re = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  sr_result_regs_r_330_Im = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  sr_result_regs_r_331_Re = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  sr_result_regs_r_331_Im = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  sr_result_regs_r_332_Re = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  sr_result_regs_r_332_Im = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  sr_result_regs_r_333_Re = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  sr_result_regs_r_333_Im = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  sr_result_regs_r_334_Re = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  sr_result_regs_r_334_Im = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  sr_result_regs_r_335_Re = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  sr_result_regs_r_335_Im = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  sr_result_regs_r_336_Re = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  sr_result_regs_r_336_Im = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  sr_result_regs_r_337_Re = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  sr_result_regs_r_337_Im = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  sr_result_regs_r_338_Re = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  sr_result_regs_r_338_Im = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  sr_result_regs_r_339_Re = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  sr_result_regs_r_339_Im = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  sr_result_regs_r_340_Re = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  sr_result_regs_r_340_Im = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  sr_result_regs_r_341_Re = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  sr_result_regs_r_341_Im = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  sr_result_regs_r_342_Re = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  sr_result_regs_r_342_Im = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  sr_result_regs_r_343_Re = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  sr_result_regs_r_343_Im = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  sr_result_regs_r_344_Re = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  sr_result_regs_r_344_Im = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  sr_result_regs_r_345_Re = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  sr_result_regs_r_345_Im = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  sr_result_regs_r_346_Re = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  sr_result_regs_r_346_Im = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  sr_result_regs_r_347_Re = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  sr_result_regs_r_347_Im = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  sr_result_regs_r_348_Re = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  sr_result_regs_r_348_Im = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  sr_result_regs_r_349_Re = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  sr_result_regs_r_349_Im = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  sr_result_regs_r_350_Re = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  sr_result_regs_r_350_Im = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  sr_result_regs_r_351_Re = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  sr_result_regs_r_351_Im = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  sr_result_regs_r_352_Re = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  sr_result_regs_r_352_Im = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  sr_result_regs_r_353_Re = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  sr_result_regs_r_353_Im = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  sr_result_regs_r_354_Re = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  sr_result_regs_r_354_Im = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  sr_result_regs_r_355_Re = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  sr_result_regs_r_355_Im = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  sr_result_regs_r_356_Re = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  sr_result_regs_r_356_Im = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  sr_result_regs_r_357_Re = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  sr_result_regs_r_357_Im = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  sr_result_regs_r_358_Re = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  sr_result_regs_r_358_Im = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  sr_result_regs_r_359_Re = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  sr_result_regs_r_359_Im = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  sr_result_regs_r_360_Re = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  sr_result_regs_r_360_Im = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  sr_result_regs_r_361_Re = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  sr_result_regs_r_361_Im = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  sr_result_regs_r_362_Re = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  sr_result_regs_r_362_Im = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  sr_result_regs_r_363_Re = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  sr_result_regs_r_363_Im = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  sr_result_regs_r_364_Re = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  sr_result_regs_r_364_Im = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  sr_result_regs_r_365_Re = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  sr_result_regs_r_365_Im = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  sr_result_regs_r_366_Re = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  sr_result_regs_r_366_Im = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  sr_result_regs_r_367_Re = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  sr_result_regs_r_367_Im = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  sr_result_regs_r_368_Re = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  sr_result_regs_r_368_Im = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  sr_result_regs_r_369_Re = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  sr_result_regs_r_369_Im = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  sr_result_regs_r_370_Re = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  sr_result_regs_r_370_Im = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  sr_result_regs_r_371_Re = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  sr_result_regs_r_371_Im = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  sr_result_regs_r_372_Re = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  sr_result_regs_r_372_Im = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  sr_result_regs_r_373_Re = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  sr_result_regs_r_373_Im = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  sr_result_regs_r_374_Re = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  sr_result_regs_r_374_Im = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  sr_result_regs_r_375_Re = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  sr_result_regs_r_375_Im = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  sr_result_regs_r_376_Re = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  sr_result_regs_r_376_Im = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  sr_result_regs_r_377_Re = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  sr_result_regs_r_377_Im = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  sr_result_regs_r_378_Re = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  sr_result_regs_r_378_Im = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  sr_result_regs_r_379_Re = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  sr_result_regs_r_379_Im = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  sr_result_regs_r_380_Re = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  sr_result_regs_r_380_Im = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  sr_result_regs_r_381_Re = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  sr_result_regs_r_381_Im = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  sr_result_regs_r_382_Re = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  sr_result_regs_r_382_Im = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  sr_result_regs_r_383_Re = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  sr_result_regs_r_383_Im = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  io_out_valid_r = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  io_out_valid_r_1 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  io_out_valid_r_2 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  io_out_valid_r_3 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  io_out_valid_r_4 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  io_out_valid_r_5 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  io_out_valid_r_6 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  io_out_valid_r_7 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  io_out_valid_r_8 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  io_out_valid_r_9 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  io_out_valid_r_10 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  io_out_valid_r_11 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  io_out_valid_r_12 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  io_out_valid_r_13 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  io_out_valid_r_14 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  io_out_valid_r_15 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  io_out_valid_r_16 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  io_out_valid_r_17 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  io_out_valid_r_18 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  io_out_valid_r_19 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  io_out_valid_r_20 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  io_out_valid_r_21 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  io_out_valid_r_22 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  io_out_valid_r_23 = _RAND_792[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32(
  input         io_in_inv,
  input  [4:0]  io_in_addr,
  output [31:0] io_out_data_0_Im,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_2_Im,
  output [31:0] io_out_data_3_Re,
  output [31:0] io_out_data_3_Im,
  output [31:0] io_out_data_4_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_6_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im,
  output [31:0] io_out_data_8_Im,
  output [31:0] io_out_data_9_Re,
  output [31:0] io_out_data_9_Im,
  output [31:0] io_out_data_10_Im,
  output [31:0] io_out_data_11_Re,
  output [31:0] io_out_data_11_Im,
  output [31:0] io_out_data_12_Im,
  output [31:0] io_out_data_13_Re,
  output [31:0] io_out_data_13_Im,
  output [31:0] io_out_data_14_Im,
  output [31:0] io_out_data_15_Re,
  output [31:0] io_out_data_15_Im
);
  wire [31:0] _GEN_10 = io_in_addr[0] ? 32'hbe14fdf0 : 32'h3f800000; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_11 = io_in_addr[0] ? 32'h3f7d4694 : 32'h0; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_14 = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_15 = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_74 = io_in_addr[0] ? 32'h3f5806d0 : 32'hbf275530; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_75 = io_in_addr[0] ? 32'hbf095cd6 : 32'hbf41bdce; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_78 = io_in_addr[0] ? 32'hbf3504f2 : 32'h3f3504f2; // @[TwidFactorDesigns.scala 26:{53,53}]
  assign io_out_data_0_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_1_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_1_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_2_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_3_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_3_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_4_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_5_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_5_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_6_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_7_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_7_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_8_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_9_Re = io_in_inv ? _GEN_74 : _GEN_78; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_9_Im = io_in_inv ? _GEN_75 : 32'hbf3504f2; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_10_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_11_Re = io_in_inv ? _GEN_74 : _GEN_78; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_11_Im = io_in_inv ? _GEN_75 : 32'hbf3504f2; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_12_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_13_Re = io_in_inv ? _GEN_74 : _GEN_78; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_13_Im = io_in_inv ? _GEN_75 : 32'hbf3504f2; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_14_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_15_Re = io_in_inv ? _GEN_74 : _GEN_78; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_15_Im = io_in_inv ? _GEN_75 : 32'hbf3504f2; // @[TwidFactorDesigns.scala 26:53]
endmodule
module multiplier_bw24(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [47:0] io_out_s
);
  assign io_out_s = io_in_a * io_in_b; // @[Arithmetic.scala 55:23]
endmodule
module twoscomplement_bw8(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _x_T = ~io_in; // @[Arithmetic.scala 13:16]
  assign io_out = 8'h1 + _x_T; // @[Arithmetic.scala 13:14]
endmodule
module full_adder_bw8(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a + io_in_b; // @[Arithmetic.scala 27:23]
  wire [9:0] _result_T_1 = {{1'd0}, _result_T}; // @[Arithmetic.scala 27:34]
  wire [8:0] result = _result_T_1[8:0]; // @[Arithmetic.scala 26:22 27:12]
  assign io_out_s = result[7:0]; // @[Arithmetic.scala 28:23]
  assign io_out_c = result[8]; // @[Arithmetic.scala 29:23]
endmodule
module FP_multiplier_bw32(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
`endif // RANDOMIZE_REG_INIT
  wire [23:0] frac_multiplier_io_in_a; // @[FPArithmetic.scala 334:33]
  wire [23:0] frac_multiplier_io_in_b; // @[FPArithmetic.scala 334:33]
  wire [47:0] frac_multiplier_io_out_s; // @[FPArithmetic.scala 334:33]
  wire [7:0] postProcess_exp_subtractor_io_in_a; // @[FPArithmetic.scala 341:44]
  wire [7:0] postProcess_exp_subtractor_io_in_b; // @[FPArithmetic.scala 341:44]
  wire [7:0] postProcess_exp_subtractor_io_out_s; // @[FPArithmetic.scala 341:44]
  wire  postProcess_exp_subtractor_io_out_c; // @[FPArithmetic.scala 341:44]
  wire [7:0] postProcess_cmpl_io_in; // @[FPArithmetic.scala 350:34]
  wire [7:0] postProcess_cmpl_io_out; // @[FPArithmetic.scala 350:34]
  wire [7:0] postProcess_exp_adder_io_in_a; // @[FPArithmetic.scala 367:39]
  wire [7:0] postProcess_exp_adder_io_in_b; // @[FPArithmetic.scala 367:39]
  wire [7:0] postProcess_exp_adder_io_out_s; // @[FPArithmetic.scala 367:39]
  wire  postProcess_exp_adder_io_out_c; // @[FPArithmetic.scala 367:39]
  wire  sign_wire_0 = io_in_a[31]; // @[FPArithmetic.scala 300:28]
  wire  sign_wire_1 = io_in_b[31]; // @[FPArithmetic.scala 301:28]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 305:64]
  wire [8:0] _GEN_62 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 305:36]
  wire [7:0] _GEN_0 = io_in_a[30:23] < 8'h1 ? 8'h1 : io_in_a[30:23]; // @[FPArithmetic.scala 307:45 308:19 310:19]
  wire [8:0] _GEN_1 = _GEN_62 > _T_2 ? _T_2 : {{1'd0}, _GEN_0}; // @[FPArithmetic.scala 305:71 306:19]
  wire [8:0] _GEN_63 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 312:36]
  wire [7:0] _GEN_2 = io_in_b[30:23] < 8'h1 ? 8'h1 : io_in_b[30:23]; // @[FPArithmetic.scala 314:45 315:19 317:19]
  wire [8:0] _GEN_3 = _GEN_63 > _T_2 ? _T_2 : {{1'd0}, _GEN_2}; // @[FPArithmetic.scala 312:71 313:19]
  wire [22:0] frac_wire_0 = io_in_a[22:0]; // @[FPArithmetic.scala 322:28]
  wire [22:0] frac_wire_1 = io_in_b[22:0]; // @[FPArithmetic.scala 323:28]
  wire [23:0] whole_frac_wire_0 = {1'h1,frac_wire_0}; // @[FPArithmetic.scala 327:31]
  wire [23:0] whole_frac_wire_1 = {1'h1,frac_wire_1}; // @[FPArithmetic.scala 328:31]
  reg  sign_reg_0_0; // @[FPArithmetic.scala 330:27]
  reg  sign_reg_0_1; // @[FPArithmetic.scala 330:27]
  reg  sign_reg_1_0; // @[FPArithmetic.scala 330:27]
  reg  sign_reg_1_1; // @[FPArithmetic.scala 330:27]
  reg  sign_reg_2_0; // @[FPArithmetic.scala 330:27]
  reg  sign_reg_2_1; // @[FPArithmetic.scala 330:27]
  reg  sign_reg_3_0; // @[FPArithmetic.scala 330:27]
  reg  sign_reg_3_1; // @[FPArithmetic.scala 330:27]
  reg  sign_reg_4_0; // @[FPArithmetic.scala 330:27]
  reg  sign_reg_4_1; // @[FPArithmetic.scala 330:27]
  reg [7:0] exp_reg_0_0; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_0_1; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_1_0; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_1_1; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_2_0; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_2_1; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_3_0; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_3_1; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_4_0; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_4_1; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_5_0; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_5_1; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_6_0; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_6_1; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_7_0; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_7_1; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_8_0; // @[FPArithmetic.scala 331:26]
  reg [7:0] exp_reg_8_1; // @[FPArithmetic.scala 331:26]
  reg [23:0] whole_frac_reg_0_0; // @[FPArithmetic.scala 332:33]
  reg [23:0] whole_frac_reg_0_1; // @[FPArithmetic.scala 332:33]
  reg [23:0] whole_frac_reg_1_0; // @[FPArithmetic.scala 332:33]
  reg [23:0] whole_frac_reg_1_1; // @[FPArithmetic.scala 332:33]
  reg [47:0] frac_multiplier_out_reg_0; // @[FPArithmetic.scala 338:42]
  reg [47:0] frac_multiplier_out_reg_1; // @[FPArithmetic.scala 338:42]
  reg [47:0] frac_multiplier_out_reg_2; // @[FPArithmetic.scala 338:42]
  reg [47:0] frac_multiplier_out_reg_3; // @[FPArithmetic.scala 338:42]
  reg [47:0] frac_multiplier_out_reg_4; // @[FPArithmetic.scala 338:42]
  reg [47:0] frac_multiplier_out_reg_5; // @[FPArithmetic.scala 338:42]
  reg [7:0] postProcess_exp_sub_out_sum_reg_0; // @[FPArithmetic.scala 346:50]
  reg [7:0] postProcess_cmpl_out_reg_0; // @[FPArithmetic.scala 353:43]
  reg [7:0] postProcess_cmpl_out_reg_1; // @[FPArithmetic.scala 353:43]
  reg [7:0] postProcess_cmpl_out_reg_2; // @[FPArithmetic.scala 353:43]
  wire  new_sign_wire = sign_reg_4_0 ^ sign_reg_4_1; // @[FPArithmetic.scala 356:37]
  reg  new_sign_reg_0; // @[FPArithmetic.scala 358:31]
  reg  new_sign_reg_1; // @[FPArithmetic.scala 358:31]
  reg  new_sign_reg_2; // @[FPArithmetic.scala 358:31]
  reg  new_sign_reg_3; // @[FPArithmetic.scala 358:31]
  wire  postProcessInstruction_wire = exp_reg_5_1 < 8'h7f; // @[FPArithmetic.scala 361:51]
  reg  postProcessInstruction_reg_0; // @[FPArithmetic.scala 363:45]
  reg  postProcessInstruction_reg_1; // @[FPArithmetic.scala 363:45]
  wire [7:0] _postProcess_exp_adder_io_in_a_T_1 = exp_reg_6_0 + 8'h1; // @[FPArithmetic.scala 371:54]
  reg [7:0] postProcess_exp_adder_out_sum_reg_0; // @[FPArithmetic.scala 378:52]
  reg  postProcess_exp_adder_out_carry_reg_0; // @[FPArithmetic.scala 379:54]
  reg [7:0] new_exp_reg_0; // @[FPArithmetic.scala 381:30]
  reg [22:0] new_frac_reg_0; // @[FPArithmetic.scala 382:31]
  reg [31:0] output_result_reg; // @[FPArithmetic.scala 384:36]
  wire  _new_exp_reg_0_T_1 = ~postProcess_exp_adder_out_carry_reg_0; // @[FPArithmetic.scala 387:64]
  wire  _new_exp_reg_0_T_5 = postProcess_exp_adder_out_carry_reg_0 | postProcess_exp_adder_out_sum_reg_0 > 8'hfe; // @[FPArithmetic.scala 387:206]
  wire [22:0] _new_frac_reg_0_T_3 = _new_exp_reg_0_T_1 ? 23'h0 : frac_multiplier_out_reg_5[46:24]; // @[FPArithmetic.scala 389:66]
  wire [22:0] _new_frac_reg_0_T_8 = _new_exp_reg_0_T_5 ? 23'h7fffff : frac_multiplier_out_reg_5[46:24]; // @[FPArithmetic.scala 389:192]
  wire [22:0] _new_frac_reg_0_T_13 = _new_exp_reg_0_T_1 ? 23'h0 : frac_multiplier_out_reg_5[45:23]; // @[FPArithmetic.scala 391:66]
  wire [22:0] _new_frac_reg_0_T_18 = _new_exp_reg_0_T_5 ? 23'h7fffff : frac_multiplier_out_reg_5[45:23]; // @[FPArithmetic.scala 391:188]
  wire [31:0] _output_result_reg_T_1 = {new_sign_reg_3,new_exp_reg_0,new_frac_reg_0}; // @[FPArithmetic.scala 426:64]
  wire [7:0] exp_wire_0 = _GEN_1[7:0]; // @[FPArithmetic.scala 304:24]
  wire [7:0] exp_wire_1 = _GEN_3[7:0]; // @[FPArithmetic.scala 304:24]
  multiplier_bw24 frac_multiplier ( // @[FPArithmetic.scala 334:33]
    .io_in_a(frac_multiplier_io_in_a),
    .io_in_b(frac_multiplier_io_in_b),
    .io_out_s(frac_multiplier_io_out_s)
  );
  full_subtractor_bw8 postProcess_exp_subtractor ( // @[FPArithmetic.scala 341:44]
    .io_in_a(postProcess_exp_subtractor_io_in_a),
    .io_in_b(postProcess_exp_subtractor_io_in_b),
    .io_out_s(postProcess_exp_subtractor_io_out_s),
    .io_out_c(postProcess_exp_subtractor_io_out_c)
  );
  twoscomplement_bw8 postProcess_cmpl ( // @[FPArithmetic.scala 350:34]
    .io_in(postProcess_cmpl_io_in),
    .io_out(postProcess_cmpl_io_out)
  );
  full_adder_bw8 postProcess_exp_adder ( // @[FPArithmetic.scala 367:39]
    .io_in_a(postProcess_exp_adder_io_in_a),
    .io_in_b(postProcess_exp_adder_io_in_b),
    .io_out_s(postProcess_exp_adder_io_out_s),
    .io_out_c(postProcess_exp_adder_io_out_c)
  );
  assign io_out_s = output_result_reg; // @[FPArithmetic.scala 429:14]
  assign frac_multiplier_io_in_a = whole_frac_reg_1_0; // @[FPArithmetic.scala 335:29]
  assign frac_multiplier_io_in_b = whole_frac_reg_1_1; // @[FPArithmetic.scala 336:29]
  assign postProcess_exp_subtractor_io_in_a = 8'h7f; // @[FPArithmetic.scala 342:40]
  assign postProcess_exp_subtractor_io_in_b = exp_reg_2_1; // @[FPArithmetic.scala 343:40]
  assign postProcess_cmpl_io_in = postProcess_exp_sub_out_sum_reg_0; // @[FPArithmetic.scala 351:28]
  assign postProcess_exp_adder_io_in_a = frac_multiplier_out_reg_4[47] ? _postProcess_exp_adder_io_in_a_T_1 :
    exp_reg_6_0; // @[FPArithmetic.scala 370:72 371:37 374:37]
  assign postProcess_exp_adder_io_in_b = postProcess_cmpl_out_reg_2; // @[FPArithmetic.scala 370:72 372:37 375:37]
  always @(posedge clock) begin
    if (reset) begin // @[FPArithmetic.scala 330:27]
      sign_reg_0_0 <= 1'h0; // @[FPArithmetic.scala 330:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      sign_reg_0_0 <= sign_wire_0; // @[FPArithmetic.scala 393:19]
    end
    if (reset) begin // @[FPArithmetic.scala 330:27]
      sign_reg_0_1 <= 1'h0; // @[FPArithmetic.scala 330:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      sign_reg_0_1 <= sign_wire_1; // @[FPArithmetic.scala 393:19]
    end
    if (reset) begin // @[FPArithmetic.scala 330:27]
      sign_reg_1_0 <= 1'h0; // @[FPArithmetic.scala 330:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      sign_reg_1_0 <= sign_reg_0_0; // @[FPArithmetic.scala 409:25]
    end
    if (reset) begin // @[FPArithmetic.scala 330:27]
      sign_reg_1_1 <= 1'h0; // @[FPArithmetic.scala 330:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      sign_reg_1_1 <= sign_reg_0_1; // @[FPArithmetic.scala 409:25]
    end
    if (reset) begin // @[FPArithmetic.scala 330:27]
      sign_reg_2_0 <= 1'h0; // @[FPArithmetic.scala 330:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      sign_reg_2_0 <= sign_reg_1_0; // @[FPArithmetic.scala 409:25]
    end
    if (reset) begin // @[FPArithmetic.scala 330:27]
      sign_reg_2_1 <= 1'h0; // @[FPArithmetic.scala 330:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      sign_reg_2_1 <= sign_reg_1_1; // @[FPArithmetic.scala 409:25]
    end
    if (reset) begin // @[FPArithmetic.scala 330:27]
      sign_reg_3_0 <= 1'h0; // @[FPArithmetic.scala 330:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      sign_reg_3_0 <= sign_reg_2_0; // @[FPArithmetic.scala 409:25]
    end
    if (reset) begin // @[FPArithmetic.scala 330:27]
      sign_reg_3_1 <= 1'h0; // @[FPArithmetic.scala 330:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      sign_reg_3_1 <= sign_reg_2_1; // @[FPArithmetic.scala 409:25]
    end
    if (reset) begin // @[FPArithmetic.scala 330:27]
      sign_reg_4_0 <= 1'h0; // @[FPArithmetic.scala 330:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      sign_reg_4_0 <= sign_reg_3_0; // @[FPArithmetic.scala 409:25]
    end
    if (reset) begin // @[FPArithmetic.scala 330:27]
      sign_reg_4_1 <= 1'h0; // @[FPArithmetic.scala 330:27]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      sign_reg_4_1 <= sign_reg_3_1; // @[FPArithmetic.scala 409:25]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_0_0 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_0_0 <= exp_wire_0; // @[FPArithmetic.scala 394:18]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_0_1 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_0_1 <= exp_wire_1; // @[FPArithmetic.scala 394:18]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_1_0 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_1_0 <= exp_reg_0_0; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_1_1 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_1_1 <= exp_reg_0_1; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_2_0 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_2_0 <= exp_reg_1_0; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_2_1 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_2_1 <= exp_reg_1_1; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_3_0 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_3_0 <= exp_reg_2_0; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_3_1 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_3_1 <= exp_reg_2_1; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_4_0 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_4_0 <= exp_reg_3_0; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_4_1 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_4_1 <= exp_reg_3_1; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_5_0 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_5_0 <= exp_reg_4_0; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_5_1 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_5_1 <= exp_reg_4_1; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_6_0 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_6_0 <= exp_reg_5_0; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_6_1 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_6_1 <= exp_reg_5_1; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_7_0 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_7_0 <= exp_reg_6_0; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_7_1 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_7_1 <= exp_reg_6_1; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_8_0 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_8_0 <= exp_reg_7_0; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 331:26]
      exp_reg_8_1 <= 8'h0; // @[FPArithmetic.scala 331:26]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      exp_reg_8_1 <= exp_reg_7_1; // @[FPArithmetic.scala 405:20]
    end
    if (reset) begin // @[FPArithmetic.scala 332:33]
      whole_frac_reg_0_0 <= 24'h0; // @[FPArithmetic.scala 332:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      whole_frac_reg_0_0 <= whole_frac_wire_0; // @[FPArithmetic.scala 395:25]
    end
    if (reset) begin // @[FPArithmetic.scala 332:33]
      whole_frac_reg_0_1 <= 24'h0; // @[FPArithmetic.scala 332:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      whole_frac_reg_0_1 <= whole_frac_wire_1; // @[FPArithmetic.scala 395:25]
    end
    if (reset) begin // @[FPArithmetic.scala 332:33]
      whole_frac_reg_1_0 <= 24'h0; // @[FPArithmetic.scala 332:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      whole_frac_reg_1_0 <= whole_frac_reg_0_0; // @[FPArithmetic.scala 415:37]
    end
    if (reset) begin // @[FPArithmetic.scala 332:33]
      whole_frac_reg_1_1 <= 24'h0; // @[FPArithmetic.scala 332:33]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      whole_frac_reg_1_1 <= whole_frac_reg_0_1; // @[FPArithmetic.scala 415:37]
    end
    if (reset) begin // @[FPArithmetic.scala 338:42]
      frac_multiplier_out_reg_0 <= 48'h0; // @[FPArithmetic.scala 338:42]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      frac_multiplier_out_reg_0 <= frac_multiplier_io_out_s; // @[FPArithmetic.scala 396:34]
    end
    if (reset) begin // @[FPArithmetic.scala 338:42]
      frac_multiplier_out_reg_1 <= 48'h0; // @[FPArithmetic.scala 338:42]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      frac_multiplier_out_reg_1 <= frac_multiplier_out_reg_0; // @[FPArithmetic.scala 407:38]
    end
    if (reset) begin // @[FPArithmetic.scala 338:42]
      frac_multiplier_out_reg_2 <= 48'h0; // @[FPArithmetic.scala 338:42]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      frac_multiplier_out_reg_2 <= frac_multiplier_out_reg_1; // @[FPArithmetic.scala 407:38]
    end
    if (reset) begin // @[FPArithmetic.scala 338:42]
      frac_multiplier_out_reg_3 <= 48'h0; // @[FPArithmetic.scala 338:42]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      frac_multiplier_out_reg_3 <= frac_multiplier_out_reg_2; // @[FPArithmetic.scala 407:38]
    end
    if (reset) begin // @[FPArithmetic.scala 338:42]
      frac_multiplier_out_reg_4 <= 48'h0; // @[FPArithmetic.scala 338:42]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      frac_multiplier_out_reg_4 <= frac_multiplier_out_reg_3; // @[FPArithmetic.scala 407:38]
    end
    if (reset) begin // @[FPArithmetic.scala 338:42]
      frac_multiplier_out_reg_5 <= 48'h0; // @[FPArithmetic.scala 338:42]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      frac_multiplier_out_reg_5 <= frac_multiplier_out_reg_4; // @[FPArithmetic.scala 407:38]
    end
    if (reset) begin // @[FPArithmetic.scala 346:50]
      postProcess_exp_sub_out_sum_reg_0 <= 8'h0; // @[FPArithmetic.scala 346:50]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      postProcess_exp_sub_out_sum_reg_0 <= postProcess_exp_subtractor_io_out_s; // @[FPArithmetic.scala 397:42]
    end
    if (reset) begin // @[FPArithmetic.scala 353:43]
      postProcess_cmpl_out_reg_0 <= 8'h0; // @[FPArithmetic.scala 353:43]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      postProcess_cmpl_out_reg_0 <= postProcess_cmpl_io_out; // @[FPArithmetic.scala 399:35]
    end
    if (reset) begin // @[FPArithmetic.scala 353:43]
      postProcess_cmpl_out_reg_1 <= 8'h0; // @[FPArithmetic.scala 353:43]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      postProcess_cmpl_out_reg_1 <= postProcess_cmpl_out_reg_0; // @[FPArithmetic.scala 413:45]
    end
    if (reset) begin // @[FPArithmetic.scala 353:43]
      postProcess_cmpl_out_reg_2 <= 8'h0; // @[FPArithmetic.scala 353:43]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      postProcess_cmpl_out_reg_2 <= postProcess_cmpl_out_reg_1; // @[FPArithmetic.scala 413:45]
    end
    if (reset) begin // @[FPArithmetic.scala 358:31]
      new_sign_reg_0 <= 1'h0; // @[FPArithmetic.scala 358:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      new_sign_reg_0 <= new_sign_wire; // @[FPArithmetic.scala 400:23]
    end
    if (reset) begin // @[FPArithmetic.scala 358:31]
      new_sign_reg_1 <= 1'h0; // @[FPArithmetic.scala 358:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      new_sign_reg_1 <= new_sign_reg_0; // @[FPArithmetic.scala 411:31]
    end
    if (reset) begin // @[FPArithmetic.scala 358:31]
      new_sign_reg_2 <= 1'h0; // @[FPArithmetic.scala 358:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      new_sign_reg_2 <= new_sign_reg_1; // @[FPArithmetic.scala 411:31]
    end
    if (reset) begin // @[FPArithmetic.scala 358:31]
      new_sign_reg_3 <= 1'h0; // @[FPArithmetic.scala 358:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      new_sign_reg_3 <= new_sign_reg_2; // @[FPArithmetic.scala 411:31]
    end
    if (reset) begin // @[FPArithmetic.scala 363:45]
      postProcessInstruction_reg_0 <= 1'h0; // @[FPArithmetic.scala 363:45]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      postProcessInstruction_reg_0 <= postProcessInstruction_wire; // @[FPArithmetic.scala 401:37]
    end
    if (reset) begin // @[FPArithmetic.scala 363:45]
      postProcessInstruction_reg_1 <= 1'h0; // @[FPArithmetic.scala 363:45]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      postProcessInstruction_reg_1 <= postProcessInstruction_reg_0; // @[FPArithmetic.scala 416:49]
    end
    if (reset) begin // @[FPArithmetic.scala 378:52]
      postProcess_exp_adder_out_sum_reg_0 <= 8'h0; // @[FPArithmetic.scala 378:52]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      postProcess_exp_adder_out_sum_reg_0 <= postProcess_exp_adder_io_out_s; // @[FPArithmetic.scala 402:44]
    end
    if (reset) begin // @[FPArithmetic.scala 379:54]
      postProcess_exp_adder_out_carry_reg_0 <= 1'h0; // @[FPArithmetic.scala 379:54]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      postProcess_exp_adder_out_carry_reg_0 <= postProcess_exp_adder_io_out_c; // @[FPArithmetic.scala 403:46]
    end
    if (reset) begin // @[FPArithmetic.scala 381:30]
      new_exp_reg_0 <= 8'h0; // @[FPArithmetic.scala 381:30]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      if (postProcessInstruction_reg_1) begin // @[FPArithmetic.scala 387:28]
        if (~postProcess_exp_adder_out_carry_reg_0) begin // @[FPArithmetic.scala 387:63]
          new_exp_reg_0 <= 8'h1;
        end else begin
          new_exp_reg_0 <= postProcess_exp_adder_out_sum_reg_0;
        end
      end else if (postProcess_exp_adder_out_carry_reg_0 | postProcess_exp_adder_out_sum_reg_0 > 8'hfe) begin // @[FPArithmetic.scala 387:159]
        new_exp_reg_0 <= 8'hfe;
      end else begin
        new_exp_reg_0 <= postProcess_exp_adder_out_sum_reg_0;
      end
    end
    if (reset) begin // @[FPArithmetic.scala 382:31]
      new_frac_reg_0 <= 23'h0; // @[FPArithmetic.scala 382:31]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      if (frac_multiplier_out_reg_5[47]) begin // @[FPArithmetic.scala 388:74]
        if (postProcessInstruction_reg_1) begin // @[FPArithmetic.scala 389:31]
          new_frac_reg_0 <= _new_frac_reg_0_T_3;
        end else begin
          new_frac_reg_0 <= _new_frac_reg_0_T_8;
        end
      end else if (postProcessInstruction_reg_1) begin // @[FPArithmetic.scala 391:31]
        new_frac_reg_0 <= _new_frac_reg_0_T_13;
      end else begin
        new_frac_reg_0 <= _new_frac_reg_0_T_18;
      end
    end
    if (reset) begin // @[FPArithmetic.scala 384:36]
      output_result_reg <= 32'h0; // @[FPArithmetic.scala 384:36]
    end else if (io_in_en) begin // @[FPArithmetic.scala 386:19]
      if (exp_reg_8_0 == 8'h0 | exp_reg_8_1 == 8'h0) begin // @[FPArithmetic.scala 423:60]
        output_result_reg <= 32'h0; // @[FPArithmetic.scala 424:27]
      end else begin
        output_result_reg <= _output_result_reg_T_1; // @[FPArithmetic.scala 426:27]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sign_reg_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sign_reg_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sign_reg_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  sign_reg_1_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  sign_reg_2_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  sign_reg_2_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  sign_reg_3_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sign_reg_3_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sign_reg_4_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sign_reg_4_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  exp_reg_0_0 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  exp_reg_0_1 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  exp_reg_1_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  exp_reg_1_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  exp_reg_2_0 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  exp_reg_2_1 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  exp_reg_3_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  exp_reg_3_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  exp_reg_4_0 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  exp_reg_4_1 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  exp_reg_5_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  exp_reg_5_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  exp_reg_6_0 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  exp_reg_6_1 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  exp_reg_7_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  exp_reg_7_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  exp_reg_8_0 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  exp_reg_8_1 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  whole_frac_reg_0_0 = _RAND_28[23:0];
  _RAND_29 = {1{`RANDOM}};
  whole_frac_reg_0_1 = _RAND_29[23:0];
  _RAND_30 = {1{`RANDOM}};
  whole_frac_reg_1_0 = _RAND_30[23:0];
  _RAND_31 = {1{`RANDOM}};
  whole_frac_reg_1_1 = _RAND_31[23:0];
  _RAND_32 = {2{`RANDOM}};
  frac_multiplier_out_reg_0 = _RAND_32[47:0];
  _RAND_33 = {2{`RANDOM}};
  frac_multiplier_out_reg_1 = _RAND_33[47:0];
  _RAND_34 = {2{`RANDOM}};
  frac_multiplier_out_reg_2 = _RAND_34[47:0];
  _RAND_35 = {2{`RANDOM}};
  frac_multiplier_out_reg_3 = _RAND_35[47:0];
  _RAND_36 = {2{`RANDOM}};
  frac_multiplier_out_reg_4 = _RAND_36[47:0];
  _RAND_37 = {2{`RANDOM}};
  frac_multiplier_out_reg_5 = _RAND_37[47:0];
  _RAND_38 = {1{`RANDOM}};
  postProcess_exp_sub_out_sum_reg_0 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  postProcess_cmpl_out_reg_0 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  postProcess_cmpl_out_reg_1 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  postProcess_cmpl_out_reg_2 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  new_sign_reg_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  new_sign_reg_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  new_sign_reg_2 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  new_sign_reg_3 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  postProcessInstruction_reg_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  postProcessInstruction_reg_1 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  postProcess_exp_adder_out_sum_reg_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  postProcess_exp_adder_out_carry_reg_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  new_exp_reg_0 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  new_frac_reg_0 = _RAND_51[22:0];
  _RAND_52 = {1{`RANDOM}};
  output_result_reg = _RAND_52[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexMultiplier_bw32(
  input         clock,
  input         reset,
  input         io_in_en,
  input         io_in_valid,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im,
  output        io_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire  FP_subtractor_bw32_clock; // @[FPComplex.scala 128:24]
  wire  FP_subtractor_bw32_reset; // @[FPComplex.scala 128:24]
  wire  FP_subtractor_bw32_io_in_en; // @[FPComplex.scala 128:24]
  wire [31:0] FP_subtractor_bw32_io_in_a; // @[FPComplex.scala 128:24]
  wire [31:0] FP_subtractor_bw32_io_in_b; // @[FPComplex.scala 128:24]
  wire [31:0] FP_subtractor_bw32_io_out_s; // @[FPComplex.scala 128:24]
  wire  FP_adder_bw32_clock; // @[FPComplex.scala 129:24]
  wire  FP_adder_bw32_reset; // @[FPComplex.scala 129:24]
  wire  FP_adder_bw32_io_in_en; // @[FPComplex.scala 129:24]
  wire [31:0] FP_adder_bw32_io_in_a; // @[FPComplex.scala 129:24]
  wire [31:0] FP_adder_bw32_io_in_b; // @[FPComplex.scala 129:24]
  wire [31:0] FP_adder_bw32_io_out_s; // @[FPComplex.scala 129:24]
  wire  FP_multiplier_bw32_clock; // @[FPComplex.scala 130:47]
  wire  FP_multiplier_bw32_reset; // @[FPComplex.scala 130:47]
  wire  FP_multiplier_bw32_io_in_en; // @[FPComplex.scala 130:47]
  wire [31:0] FP_multiplier_bw32_io_in_a; // @[FPComplex.scala 130:47]
  wire [31:0] FP_multiplier_bw32_io_in_b; // @[FPComplex.scala 130:47]
  wire [31:0] FP_multiplier_bw32_io_out_s; // @[FPComplex.scala 130:47]
  wire  FP_multiplier_bw32_1_clock; // @[FPComplex.scala 130:47]
  wire  FP_multiplier_bw32_1_reset; // @[FPComplex.scala 130:47]
  wire  FP_multiplier_bw32_1_io_in_en; // @[FPComplex.scala 130:47]
  wire [31:0] FP_multiplier_bw32_1_io_in_a; // @[FPComplex.scala 130:47]
  wire [31:0] FP_multiplier_bw32_1_io_in_b; // @[FPComplex.scala 130:47]
  wire [31:0] FP_multiplier_bw32_1_io_out_s; // @[FPComplex.scala 130:47]
  wire  FP_multiplier_bw32_2_clock; // @[FPComplex.scala 130:47]
  wire  FP_multiplier_bw32_2_reset; // @[FPComplex.scala 130:47]
  wire  FP_multiplier_bw32_2_io_in_en; // @[FPComplex.scala 130:47]
  wire [31:0] FP_multiplier_bw32_2_io_in_a; // @[FPComplex.scala 130:47]
  wire [31:0] FP_multiplier_bw32_2_io_in_b; // @[FPComplex.scala 130:47]
  wire [31:0] FP_multiplier_bw32_2_io_out_s; // @[FPComplex.scala 130:47]
  wire  FP_multiplier_bw32_3_clock; // @[FPComplex.scala 130:47]
  wire  FP_multiplier_bw32_3_reset; // @[FPComplex.scala 130:47]
  wire  FP_multiplier_bw32_3_io_in_en; // @[FPComplex.scala 130:47]
  wire [31:0] FP_multiplier_bw32_3_io_in_a; // @[FPComplex.scala 130:47]
  wire [31:0] FP_multiplier_bw32_3_io_in_b; // @[FPComplex.scala 130:47]
  wire [31:0] FP_multiplier_bw32_3_io_out_s; // @[FPComplex.scala 130:47]
  reg  io_out_valid_r; // @[Reg.scala 16:16]
  reg  io_out_valid_r_1; // @[Reg.scala 16:16]
  reg  io_out_valid_r_2; // @[Reg.scala 16:16]
  reg  io_out_valid_r_3; // @[Reg.scala 16:16]
  reg  io_out_valid_r_4; // @[Reg.scala 16:16]
  reg  io_out_valid_r_5; // @[Reg.scala 16:16]
  reg  io_out_valid_r_6; // @[Reg.scala 16:16]
  reg  io_out_valid_r_7; // @[Reg.scala 16:16]
  reg  io_out_valid_r_8; // @[Reg.scala 16:16]
  reg  io_out_valid_r_9; // @[Reg.scala 16:16]
  reg  io_out_valid_r_10; // @[Reg.scala 16:16]
  reg  io_out_valid_r_11; // @[Reg.scala 16:16]
  reg  io_out_valid_r_12; // @[Reg.scala 16:16]
  reg  io_out_valid_r_13; // @[Reg.scala 16:16]
  reg  io_out_valid_r_14; // @[Reg.scala 16:16]
  reg  io_out_valid_r_15; // @[Reg.scala 16:16]
  reg  io_out_valid_r_16; // @[Reg.scala 16:16]
  reg  io_out_valid_r_17; // @[Reg.scala 16:16]
  reg  io_out_valid_r_18; // @[Reg.scala 16:16]
  reg  io_out_valid_r_19; // @[Reg.scala 16:16]
  reg  io_out_valid_r_20; // @[Reg.scala 16:16]
  reg  io_out_valid_r_21; // @[Reg.scala 16:16]
  reg  io_out_valid_r_22; // @[Reg.scala 16:16]
  FP_subtractor_bw32 FP_subtractor_bw32 ( // @[FPComplex.scala 128:24]
    .clock(FP_subtractor_bw32_clock),
    .reset(FP_subtractor_bw32_reset),
    .io_in_en(FP_subtractor_bw32_io_in_en),
    .io_in_a(FP_subtractor_bw32_io_in_a),
    .io_in_b(FP_subtractor_bw32_io_in_b),
    .io_out_s(FP_subtractor_bw32_io_out_s)
  );
  FP_adder_bw32 FP_adder_bw32 ( // @[FPComplex.scala 129:24]
    .clock(FP_adder_bw32_clock),
    .reset(FP_adder_bw32_reset),
    .io_in_en(FP_adder_bw32_io_in_en),
    .io_in_a(FP_adder_bw32_io_in_a),
    .io_in_b(FP_adder_bw32_io_in_b),
    .io_out_s(FP_adder_bw32_io_out_s)
  );
  FP_multiplier_bw32 FP_multiplier_bw32 ( // @[FPComplex.scala 130:47]
    .clock(FP_multiplier_bw32_clock),
    .reset(FP_multiplier_bw32_reset),
    .io_in_en(FP_multiplier_bw32_io_in_en),
    .io_in_a(FP_multiplier_bw32_io_in_a),
    .io_in_b(FP_multiplier_bw32_io_in_b),
    .io_out_s(FP_multiplier_bw32_io_out_s)
  );
  FP_multiplier_bw32 FP_multiplier_bw32_1 ( // @[FPComplex.scala 130:47]
    .clock(FP_multiplier_bw32_1_clock),
    .reset(FP_multiplier_bw32_1_reset),
    .io_in_en(FP_multiplier_bw32_1_io_in_en),
    .io_in_a(FP_multiplier_bw32_1_io_in_a),
    .io_in_b(FP_multiplier_bw32_1_io_in_b),
    .io_out_s(FP_multiplier_bw32_1_io_out_s)
  );
  FP_multiplier_bw32 FP_multiplier_bw32_2 ( // @[FPComplex.scala 130:47]
    .clock(FP_multiplier_bw32_2_clock),
    .reset(FP_multiplier_bw32_2_reset),
    .io_in_en(FP_multiplier_bw32_2_io_in_en),
    .io_in_a(FP_multiplier_bw32_2_io_in_a),
    .io_in_b(FP_multiplier_bw32_2_io_in_b),
    .io_out_s(FP_multiplier_bw32_2_io_out_s)
  );
  FP_multiplier_bw32 FP_multiplier_bw32_3 ( // @[FPComplex.scala 130:47]
    .clock(FP_multiplier_bw32_3_clock),
    .reset(FP_multiplier_bw32_3_reset),
    .io_in_en(FP_multiplier_bw32_3_io_in_en),
    .io_in_a(FP_multiplier_bw32_3_io_in_a),
    .io_in_b(FP_multiplier_bw32_3_io_in_b),
    .io_out_s(FP_multiplier_bw32_3_io_out_s)
  );
  assign io_out_s_Re = FP_subtractor_bw32_io_out_s; // @[FPComplex.scala 146:17]
  assign io_out_s_Im = FP_adder_bw32_io_out_s; // @[FPComplex.scala 147:17]
  assign io_out_valid = io_out_valid_r_22; // @[FPComplex.scala 148:18]
  assign FP_subtractor_bw32_clock = clock;
  assign FP_subtractor_bw32_reset = reset;
  assign FP_subtractor_bw32_io_in_en = io_in_en; // @[FPComplex.scala 132:18]
  assign FP_subtractor_bw32_io_in_a = FP_multiplier_bw32_io_out_s; // @[FPComplex.scala 142:17]
  assign FP_subtractor_bw32_io_in_b = FP_multiplier_bw32_1_io_out_s; // @[FPComplex.scala 143:17]
  assign FP_adder_bw32_clock = clock;
  assign FP_adder_bw32_reset = reset;
  assign FP_adder_bw32_io_in_en = io_in_en; // @[FPComplex.scala 133:18]
  assign FP_adder_bw32_io_in_a = FP_multiplier_bw32_2_io_out_s; // @[FPComplex.scala 144:17]
  assign FP_adder_bw32_io_in_b = FP_multiplier_bw32_3_io_out_s; // @[FPComplex.scala 145:17]
  assign FP_multiplier_bw32_clock = clock;
  assign FP_multiplier_bw32_reset = reset;
  assign FP_multiplier_bw32_io_in_en = io_in_en; // @[FPComplex.scala 131:36]
  assign FP_multiplier_bw32_io_in_a = io_in_a_Re; // @[FPComplex.scala 134:28]
  assign FP_multiplier_bw32_io_in_b = io_in_b_Re; // @[FPComplex.scala 135:28]
  assign FP_multiplier_bw32_1_clock = clock;
  assign FP_multiplier_bw32_1_reset = reset;
  assign FP_multiplier_bw32_1_io_in_en = io_in_en; // @[FPComplex.scala 131:36]
  assign FP_multiplier_bw32_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 136:28]
  assign FP_multiplier_bw32_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 137:28]
  assign FP_multiplier_bw32_2_clock = clock;
  assign FP_multiplier_bw32_2_reset = reset;
  assign FP_multiplier_bw32_2_io_in_en = io_in_en; // @[FPComplex.scala 131:36]
  assign FP_multiplier_bw32_2_io_in_a = io_in_a_Re; // @[FPComplex.scala 138:28]
  assign FP_multiplier_bw32_2_io_in_b = io_in_b_Im; // @[FPComplex.scala 139:28]
  assign FP_multiplier_bw32_3_clock = clock;
  assign FP_multiplier_bw32_3_reset = reset;
  assign FP_multiplier_bw32_3_io_in_en = io_in_en; // @[FPComplex.scala 131:36]
  assign FP_multiplier_bw32_3_io_in_a = io_in_a_Im; // @[FPComplex.scala 140:28]
  assign FP_multiplier_bw32_3_io_in_b = io_in_b_Re; // @[FPComplex.scala 141:28]
  always @(posedge clock) begin
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r <= io_in_valid; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_1 <= io_out_valid_r; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_2 <= io_out_valid_r_1; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_3 <= io_out_valid_r_2; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_4 <= io_out_valid_r_3; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_5 <= io_out_valid_r_4; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_6 <= io_out_valid_r_5; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_7 <= io_out_valid_r_6; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_8 <= io_out_valid_r_7; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_9 <= io_out_valid_r_8; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_10 <= io_out_valid_r_9; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_11 <= io_out_valid_r_10; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_12 <= io_out_valid_r_11; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_13 <= io_out_valid_r_12; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_14 <= io_out_valid_r_13; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_15 <= io_out_valid_r_14; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_16 <= io_out_valid_r_15; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_17 <= io_out_valid_r_16; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_18 <= io_out_valid_r_17; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_19 <= io_out_valid_r_18; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_20 <= io_out_valid_r_19; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_21 <= io_out_valid_r_20; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r_22 <= io_out_valid_r_21; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_valid_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_out_valid_r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_out_valid_r_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  io_out_valid_r_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_out_valid_r_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  io_out_valid_r_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  io_out_valid_r_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_out_valid_r_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_out_valid_r_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  io_out_valid_r_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_out_valid_r_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  io_out_valid_r_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  io_out_valid_r_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  io_out_valid_r_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  io_out_valid_r_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  io_out_valid_r_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  io_out_valid_r_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  io_out_valid_r_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  io_out_valid_r_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  io_out_valid_r_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  io_out_valid_r_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  io_out_valid_r_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  io_out_valid_r_22 = _RAND_22[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32(
  input         clock,
  input         reset,
  input         io_in_inv,
  input         io_in_en,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_valid,
  output        io_out_valid,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  wire  TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_inv; // @[TwidFactorDesigns.scala 49:28]
  wire [4:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_addr; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_0_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_1_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_1_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_2_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_3_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_3_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_4_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_5_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_5_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_6_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_7_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_7_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_8_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_9_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_9_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_10_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_11_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_11_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_12_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_13_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_13_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_14_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_15_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_15_Im; // @[TwidFactorDesigns.scala 49:28]
  wire  FPComplexMultiplier_bw32_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  reg  value_1; // @[Counter.scala 62:40]
  wire  _value_T_1 = value_1 + 1'h1; // @[Counter.scala 78:24]
  reg [31:0] multipliers_sr_out_r_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_1_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_1_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_2_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_2_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_3_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_3_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_4_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_4_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_5_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_5_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_6_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_6_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_7_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_7_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_8_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_8_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_9_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_9_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_10_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_10_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_11_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_11_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_12_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_12_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_13_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_13_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_14_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_14_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_15_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_15_Im; // @[Reg.scala 16:16]
  reg  io_out_valid_r; // @[Reg.scala 16:16]
  TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32 TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32 ( // @[TwidFactorDesigns.scala 49:28]
    .io_in_inv(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_inv),
    .io_in_addr(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_addr),
    .io_out_data_0_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_0_Im),
    .io_out_data_1_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_1_Im),
    .io_out_data_2_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_2_Im),
    .io_out_data_3_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_3_Re),
    .io_out_data_3_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_3_Im),
    .io_out_data_4_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_4_Im),
    .io_out_data_5_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_5_Im),
    .io_out_data_6_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_6_Im),
    .io_out_data_7_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_7_Im),
    .io_out_data_8_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_8_Im),
    .io_out_data_9_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_9_Re),
    .io_out_data_9_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_9_Im),
    .io_out_data_10_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_10_Im),
    .io_out_data_11_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_11_Re),
    .io_out_data_11_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_11_Im),
    .io_out_data_12_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_12_Im),
    .io_out_data_13_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_13_Re),
    .io_out_data_13_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_13_Im),
    .io_out_data_14_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_14_Im),
    .io_out_data_15_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_15_Re),
    .io_out_data_15_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_15_Im)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_clock),
    .reset(FPComplexMultiplier_bw32_reset),
    .io_in_en(FPComplexMultiplier_bw32_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_1 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_1_clock),
    .reset(FPComplexMultiplier_bw32_1_reset),
    .io_in_en(FPComplexMultiplier_bw32_1_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_1_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_1_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_1_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_2 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_2_clock),
    .reset(FPComplexMultiplier_bw32_2_reset),
    .io_in_en(FPComplexMultiplier_bw32_2_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_2_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_2_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_2_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_3 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_3_clock),
    .reset(FPComplexMultiplier_bw32_3_reset),
    .io_in_en(FPComplexMultiplier_bw32_3_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_3_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_3_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_3_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_4 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_4_clock),
    .reset(FPComplexMultiplier_bw32_4_reset),
    .io_in_en(FPComplexMultiplier_bw32_4_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_4_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_4_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_4_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_5 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_5_clock),
    .reset(FPComplexMultiplier_bw32_5_reset),
    .io_in_en(FPComplexMultiplier_bw32_5_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_5_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_5_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_5_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_6 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_6_clock),
    .reset(FPComplexMultiplier_bw32_6_reset),
    .io_in_en(FPComplexMultiplier_bw32_6_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_6_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_6_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_6_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_7 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_7_clock),
    .reset(FPComplexMultiplier_bw32_7_reset),
    .io_in_en(FPComplexMultiplier_bw32_7_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_7_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_7_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_7_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_8 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_8_clock),
    .reset(FPComplexMultiplier_bw32_8_reset),
    .io_in_en(FPComplexMultiplier_bw32_8_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_8_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_8_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_8_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_8_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_8_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_8_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_9 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_9_clock),
    .reset(FPComplexMultiplier_bw32_9_reset),
    .io_in_en(FPComplexMultiplier_bw32_9_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_9_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_9_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_9_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_10 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_10_clock),
    .reset(FPComplexMultiplier_bw32_10_reset),
    .io_in_en(FPComplexMultiplier_bw32_10_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_10_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_10_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_10_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_10_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_10_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_10_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_11 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_11_clock),
    .reset(FPComplexMultiplier_bw32_11_reset),
    .io_in_en(FPComplexMultiplier_bw32_11_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_11_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_11_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_11_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_12 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_12_clock),
    .reset(FPComplexMultiplier_bw32_12_reset),
    .io_in_en(FPComplexMultiplier_bw32_12_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_12_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_12_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_12_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_12_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_12_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_12_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_13 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_13_clock),
    .reset(FPComplexMultiplier_bw32_13_reset),
    .io_in_en(FPComplexMultiplier_bw32_13_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_13_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_13_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_13_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_14 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_14_clock),
    .reset(FPComplexMultiplier_bw32_14_reset),
    .io_in_en(FPComplexMultiplier_bw32_14_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_14_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_14_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_14_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_14_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_14_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_14_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_15 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_15_clock),
    .reset(FPComplexMultiplier_bw32_15_reset),
    .io_in_en(FPComplexMultiplier_bw32_15_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_15_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_15_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_15_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_15_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_15_io_out_valid)
  );
  assign io_out_valid = io_out_valid_r; // @[TwidFactorDesigns.scala 77:22]
  assign io_out_0_Re = multipliers_sr_out_r_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_0_Im = multipliers_sr_out_r_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_1_Re = multipliers_sr_out_r_1_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_1_Im = multipliers_sr_out_r_1_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_2_Re = multipliers_sr_out_r_2_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_2_Im = multipliers_sr_out_r_2_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_3_Re = multipliers_sr_out_r_3_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_3_Im = multipliers_sr_out_r_3_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_4_Re = multipliers_sr_out_r_4_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_4_Im = multipliers_sr_out_r_4_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_5_Re = multipliers_sr_out_r_5_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_5_Im = multipliers_sr_out_r_5_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_6_Re = multipliers_sr_out_r_6_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_6_Im = multipliers_sr_out_r_6_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_7_Re = multipliers_sr_out_r_7_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_7_Im = multipliers_sr_out_r_7_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_8_Re = multipliers_sr_out_r_8_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_8_Im = multipliers_sr_out_r_8_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_9_Re = multipliers_sr_out_r_9_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_9_Im = multipliers_sr_out_r_9_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_10_Re = multipliers_sr_out_r_10_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_10_Im = multipliers_sr_out_r_10_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_11_Re = multipliers_sr_out_r_11_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_11_Im = multipliers_sr_out_r_11_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_12_Re = multipliers_sr_out_r_12_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_12_Im = multipliers_sr_out_r_12_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_13_Re = multipliers_sr_out_r_13_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_13_Im = multipliers_sr_out_r_13_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_14_Re = multipliers_sr_out_r_14_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_14_Im = multipliers_sr_out_r_14_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_15_Re = multipliers_sr_out_r_15_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_15_Im = multipliers_sr_out_r_15_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_inv = io_in_inv; // @[TwidFactorDesigns.scala 56:23]
  assign TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_addr = {{4'd0}, value_1}; // @[TwidFactorDesigns.scala 55:24]
  assign FPComplexMultiplier_bw32_clock = clock;
  assign FPComplexMultiplier_bw32_reset = reset;
  assign FPComplexMultiplier_bw32_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_io_in_a_Re = io_in_0_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_io_in_a_Im = io_in_0_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_0_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_1_clock = clock;
  assign FPComplexMultiplier_bw32_1_reset = reset;
  assign FPComplexMultiplier_bw32_1_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_1_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_1_io_in_a_Re = io_in_1_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_1_io_in_a_Im = io_in_1_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_1_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_1_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_1_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_1_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_2_clock = clock;
  assign FPComplexMultiplier_bw32_2_reset = reset;
  assign FPComplexMultiplier_bw32_2_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_2_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_2_io_in_a_Re = io_in_2_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_2_io_in_a_Im = io_in_2_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_2_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_2_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_2_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_3_clock = clock;
  assign FPComplexMultiplier_bw32_3_reset = reset;
  assign FPComplexMultiplier_bw32_3_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_3_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_3_io_in_a_Re = io_in_3_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_3_io_in_a_Im = io_in_3_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_3_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_3_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_3_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_3_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_4_clock = clock;
  assign FPComplexMultiplier_bw32_4_reset = reset;
  assign FPComplexMultiplier_bw32_4_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_4_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_4_io_in_a_Re = io_in_4_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_4_io_in_a_Im = io_in_4_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_4_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_4_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_4_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_5_clock = clock;
  assign FPComplexMultiplier_bw32_5_reset = reset;
  assign FPComplexMultiplier_bw32_5_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_5_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_5_io_in_a_Re = io_in_5_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_5_io_in_a_Im = io_in_5_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_5_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_5_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_5_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_5_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_6_clock = clock;
  assign FPComplexMultiplier_bw32_6_reset = reset;
  assign FPComplexMultiplier_bw32_6_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_6_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_6_io_in_a_Re = io_in_6_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_6_io_in_a_Im = io_in_6_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_6_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_6_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_6_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_7_clock = clock;
  assign FPComplexMultiplier_bw32_7_reset = reset;
  assign FPComplexMultiplier_bw32_7_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_7_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_7_io_in_a_Re = io_in_7_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_7_io_in_a_Im = io_in_7_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_7_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_7_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_7_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_7_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_8_clock = clock;
  assign FPComplexMultiplier_bw32_8_reset = reset;
  assign FPComplexMultiplier_bw32_8_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_8_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_8_io_in_a_Re = io_in_8_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_8_io_in_a_Im = io_in_8_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_8_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_8_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_8_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_9_clock = clock;
  assign FPComplexMultiplier_bw32_9_reset = reset;
  assign FPComplexMultiplier_bw32_9_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_9_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_9_io_in_a_Re = io_in_9_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_9_io_in_a_Im = io_in_9_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_9_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_9_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_9_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_9_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_10_clock = clock;
  assign FPComplexMultiplier_bw32_10_reset = reset;
  assign FPComplexMultiplier_bw32_10_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_10_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_10_io_in_a_Re = io_in_10_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_10_io_in_a_Im = io_in_10_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_10_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_10_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_10_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_11_clock = clock;
  assign FPComplexMultiplier_bw32_11_reset = reset;
  assign FPComplexMultiplier_bw32_11_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_11_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_11_io_in_a_Re = io_in_11_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_11_io_in_a_Im = io_in_11_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_11_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_11_Re
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_11_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_11_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_12_clock = clock;
  assign FPComplexMultiplier_bw32_12_reset = reset;
  assign FPComplexMultiplier_bw32_12_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_12_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_12_io_in_a_Re = io_in_12_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_12_io_in_a_Im = io_in_12_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_12_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_12_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_12_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_13_clock = clock;
  assign FPComplexMultiplier_bw32_13_reset = reset;
  assign FPComplexMultiplier_bw32_13_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_13_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_13_io_in_a_Re = io_in_13_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_13_io_in_a_Im = io_in_13_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_13_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_13_Re
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_13_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_13_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_14_clock = clock;
  assign FPComplexMultiplier_bw32_14_reset = reset;
  assign FPComplexMultiplier_bw32_14_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_14_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_14_io_in_a_Re = io_in_14_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_14_io_in_a_Im = io_in_14_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_14_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_14_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_14_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_15_clock = clock;
  assign FPComplexMultiplier_bw32_15_reset = reset;
  assign FPComplexMultiplier_bw32_15_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_15_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_15_io_in_a_Re = io_in_15_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_15_io_in_a_Im = io_in_15_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_15_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_15_Re
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_15_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_data_15_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en) begin // @[TwidFactorDesigns.scala 57:22]
      if (io_in_valid) begin // @[TwidFactorDesigns.scala 58:27]
        value_1 <= _value_T_1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_Re <= FPComplexMultiplier_bw32_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_Im <= FPComplexMultiplier_bw32_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_1_Re <= FPComplexMultiplier_bw32_1_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_1_Im <= FPComplexMultiplier_bw32_1_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_2_Re <= FPComplexMultiplier_bw32_2_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_2_Im <= FPComplexMultiplier_bw32_2_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_3_Re <= FPComplexMultiplier_bw32_3_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_3_Im <= FPComplexMultiplier_bw32_3_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_4_Re <= FPComplexMultiplier_bw32_4_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_4_Im <= FPComplexMultiplier_bw32_4_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_5_Re <= FPComplexMultiplier_bw32_5_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_5_Im <= FPComplexMultiplier_bw32_5_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_6_Re <= FPComplexMultiplier_bw32_6_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_6_Im <= FPComplexMultiplier_bw32_6_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_7_Re <= FPComplexMultiplier_bw32_7_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_7_Im <= FPComplexMultiplier_bw32_7_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_8_Re <= FPComplexMultiplier_bw32_8_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_8_Im <= FPComplexMultiplier_bw32_8_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_9_Re <= FPComplexMultiplier_bw32_9_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_9_Im <= FPComplexMultiplier_bw32_9_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_10_Re <= FPComplexMultiplier_bw32_10_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_10_Im <= FPComplexMultiplier_bw32_10_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_11_Re <= FPComplexMultiplier_bw32_11_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_11_Im <= FPComplexMultiplier_bw32_11_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_12_Re <= FPComplexMultiplier_bw32_12_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_12_Im <= FPComplexMultiplier_bw32_12_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_13_Re <= FPComplexMultiplier_bw32_13_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_13_Im <= FPComplexMultiplier_bw32_13_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_14_Re <= FPComplexMultiplier_bw32_14_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_14_Im <= FPComplexMultiplier_bw32_14_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_15_Re <= FPComplexMultiplier_bw32_15_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_15_Im <= FPComplexMultiplier_bw32_15_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r <= FPComplexMultiplier_bw32_io_out_valid; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  multipliers_sr_out_r_Re = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  multipliers_sr_out_r_Im = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  multipliers_sr_out_r_1_Re = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  multipliers_sr_out_r_1_Im = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  multipliers_sr_out_r_2_Re = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  multipliers_sr_out_r_2_Im = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  multipliers_sr_out_r_3_Re = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  multipliers_sr_out_r_3_Im = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  multipliers_sr_out_r_4_Re = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  multipliers_sr_out_r_4_Im = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  multipliers_sr_out_r_5_Re = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  multipliers_sr_out_r_5_Im = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  multipliers_sr_out_r_6_Re = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  multipliers_sr_out_r_6_Im = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  multipliers_sr_out_r_7_Re = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  multipliers_sr_out_r_7_Im = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  multipliers_sr_out_r_8_Re = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  multipliers_sr_out_r_8_Im = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  multipliers_sr_out_r_9_Re = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  multipliers_sr_out_r_9_Im = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  multipliers_sr_out_r_10_Re = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  multipliers_sr_out_r_10_Im = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  multipliers_sr_out_r_11_Re = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  multipliers_sr_out_r_11_Im = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  multipliers_sr_out_r_12_Re = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  multipliers_sr_out_r_12_Im = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  multipliers_sr_out_r_13_Re = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  multipliers_sr_out_r_13_Im = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  multipliers_sr_out_r_14_Re = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  multipliers_sr_out_r_14_Im = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  multipliers_sr_out_r_15_Re = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  multipliers_sr_out_r_15_Im = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  io_out_valid_r = _RAND_33[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32(
  input         io_in_inv,
  input  [4:0]  io_in_addr,
  output [31:0] io_out_data_0_Im,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_2_Im,
  output [31:0] io_out_data_3_Re,
  output [31:0] io_out_data_3_Im,
  output [31:0] io_out_data_4_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_6_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im,
  output [31:0] io_out_data_8_Im,
  output [31:0] io_out_data_9_Re,
  output [31:0] io_out_data_9_Im,
  output [31:0] io_out_data_10_Im,
  output [31:0] io_out_data_11_Re,
  output [31:0] io_out_data_11_Im,
  output [31:0] io_out_data_12_Im,
  output [31:0] io_out_data_13_Re,
  output [31:0] io_out_data_13_Im,
  output [31:0] io_out_data_14_Im,
  output [31:0] io_out_data_15_Re,
  output [31:0] io_out_data_15_Im
);
  wire [31:0] _GEN_10 = io_in_addr[0] ? 32'hbe14fdf0 : 32'h3f800000; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_11 = io_in_addr[0] ? 32'h3f7d4694 : 32'h0; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_14 = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_15 = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_42 = io_in_addr[0] ? 32'hbf56cd64 : 32'hbed51130; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_43 = io_in_addr[0] ? 32'hbf0b44f6 : 32'h3f68c7b6; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_46 = io_in_addr[0] ? 32'hbec3ef14 : 32'h3f6c835e; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_47 = io_in_addr[0] ? 32'hbf6c835e : 32'hbec3ef14; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_74 = io_in_addr[0] ? 32'h3f5806d0 : 32'hbf275530; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_75 = io_in_addr[0] ? 32'hbf095cd6 : 32'hbf41bdce; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_78 = io_in_addr[0] ? 32'hbf3504f2 : 32'h3f3504f2; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_106 = io_in_addr[0] ? 32'h3e0c04d0 : 32'h3f75cdb8; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_107 = io_in_addr[0] ? 32'h3f7d9870 : 32'hbe8f0f8c; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_110 = io_in_addr[0] ? 32'hbf6c835e : 32'h3ec3ef14; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_111 = io_in_addr[0] ? 32'hbec3ef14 : 32'hbf6c835e; // @[TwidFactorDesigns.scala 26:{53,53}]
  assign io_out_data_0_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_1_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_1_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_2_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_3_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_3_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_4_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_5_Re = io_in_inv ? _GEN_42 : _GEN_46; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_5_Im = io_in_inv ? _GEN_43 : _GEN_47; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_6_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_7_Re = io_in_inv ? _GEN_42 : _GEN_46; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_7_Im = io_in_inv ? _GEN_43 : _GEN_47; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_8_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_9_Re = io_in_inv ? _GEN_74 : _GEN_78; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_9_Im = io_in_inv ? _GEN_75 : 32'hbf3504f2; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_10_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_11_Re = io_in_inv ? _GEN_74 : _GEN_78; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_11_Im = io_in_inv ? _GEN_75 : 32'hbf3504f2; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_12_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_13_Re = io_in_inv ? _GEN_106 : _GEN_110; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_13_Im = io_in_inv ? _GEN_107 : _GEN_111; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_14_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_15_Re = io_in_inv ? _GEN_106 : _GEN_110; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_15_Im = io_in_inv ? _GEN_107 : _GEN_111; // @[TwidFactorDesigns.scala 26:53]
endmodule
module TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32(
  input         clock,
  input         reset,
  input         io_in_inv,
  input         io_in_en,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_valid,
  output        io_out_valid,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  wire  TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_inv; // @[TwidFactorDesigns.scala 49:28]
  wire [4:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_addr; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_0_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_1_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_1_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_2_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_3_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_3_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_4_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_5_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_5_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_6_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_7_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_7_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_8_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_9_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_9_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_10_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_11_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_11_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_12_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_13_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_13_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_14_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_15_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_15_Im; // @[TwidFactorDesigns.scala 49:28]
  wire  FPComplexMultiplier_bw32_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  reg  value_1; // @[Counter.scala 62:40]
  wire  _value_T_1 = value_1 + 1'h1; // @[Counter.scala 78:24]
  reg [31:0] multipliers_sr_out_r_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_1_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_1_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_2_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_2_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_3_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_3_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_4_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_4_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_5_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_5_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_6_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_6_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_7_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_7_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_8_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_8_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_9_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_9_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_10_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_10_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_11_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_11_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_12_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_12_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_13_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_13_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_14_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_14_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_15_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_15_Im; // @[Reg.scala 16:16]
  reg  io_out_valid_r; // @[Reg.scala 16:16]
  TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32 TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32 ( // @[TwidFactorDesigns.scala 49:28]
    .io_in_inv(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_inv),
    .io_in_addr(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_addr),
    .io_out_data_0_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_0_Im),
    .io_out_data_1_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_1_Im),
    .io_out_data_2_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_2_Im),
    .io_out_data_3_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_3_Re),
    .io_out_data_3_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_3_Im),
    .io_out_data_4_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_4_Im),
    .io_out_data_5_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_5_Im),
    .io_out_data_6_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_6_Im),
    .io_out_data_7_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_7_Im),
    .io_out_data_8_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_8_Im),
    .io_out_data_9_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_9_Re),
    .io_out_data_9_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_9_Im),
    .io_out_data_10_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_10_Im),
    .io_out_data_11_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_11_Re),
    .io_out_data_11_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_11_Im),
    .io_out_data_12_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_12_Im),
    .io_out_data_13_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_13_Re),
    .io_out_data_13_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_13_Im),
    .io_out_data_14_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_14_Im),
    .io_out_data_15_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_15_Re),
    .io_out_data_15_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_15_Im)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_clock),
    .reset(FPComplexMultiplier_bw32_reset),
    .io_in_en(FPComplexMultiplier_bw32_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_1 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_1_clock),
    .reset(FPComplexMultiplier_bw32_1_reset),
    .io_in_en(FPComplexMultiplier_bw32_1_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_1_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_1_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_1_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_2 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_2_clock),
    .reset(FPComplexMultiplier_bw32_2_reset),
    .io_in_en(FPComplexMultiplier_bw32_2_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_2_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_2_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_2_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_3 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_3_clock),
    .reset(FPComplexMultiplier_bw32_3_reset),
    .io_in_en(FPComplexMultiplier_bw32_3_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_3_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_3_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_3_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_4 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_4_clock),
    .reset(FPComplexMultiplier_bw32_4_reset),
    .io_in_en(FPComplexMultiplier_bw32_4_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_4_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_4_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_4_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_5 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_5_clock),
    .reset(FPComplexMultiplier_bw32_5_reset),
    .io_in_en(FPComplexMultiplier_bw32_5_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_5_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_5_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_5_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_6 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_6_clock),
    .reset(FPComplexMultiplier_bw32_6_reset),
    .io_in_en(FPComplexMultiplier_bw32_6_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_6_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_6_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_6_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_7 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_7_clock),
    .reset(FPComplexMultiplier_bw32_7_reset),
    .io_in_en(FPComplexMultiplier_bw32_7_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_7_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_7_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_7_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_8 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_8_clock),
    .reset(FPComplexMultiplier_bw32_8_reset),
    .io_in_en(FPComplexMultiplier_bw32_8_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_8_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_8_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_8_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_8_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_8_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_8_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_9 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_9_clock),
    .reset(FPComplexMultiplier_bw32_9_reset),
    .io_in_en(FPComplexMultiplier_bw32_9_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_9_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_9_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_9_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_10 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_10_clock),
    .reset(FPComplexMultiplier_bw32_10_reset),
    .io_in_en(FPComplexMultiplier_bw32_10_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_10_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_10_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_10_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_10_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_10_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_10_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_11 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_11_clock),
    .reset(FPComplexMultiplier_bw32_11_reset),
    .io_in_en(FPComplexMultiplier_bw32_11_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_11_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_11_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_11_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_12 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_12_clock),
    .reset(FPComplexMultiplier_bw32_12_reset),
    .io_in_en(FPComplexMultiplier_bw32_12_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_12_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_12_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_12_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_12_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_12_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_12_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_13 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_13_clock),
    .reset(FPComplexMultiplier_bw32_13_reset),
    .io_in_en(FPComplexMultiplier_bw32_13_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_13_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_13_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_13_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_14 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_14_clock),
    .reset(FPComplexMultiplier_bw32_14_reset),
    .io_in_en(FPComplexMultiplier_bw32_14_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_14_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_14_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_14_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_14_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_14_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_14_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_15 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_15_clock),
    .reset(FPComplexMultiplier_bw32_15_reset),
    .io_in_en(FPComplexMultiplier_bw32_15_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_15_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_15_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_15_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_15_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_15_io_out_valid)
  );
  assign io_out_valid = io_out_valid_r; // @[TwidFactorDesigns.scala 77:22]
  assign io_out_0_Re = multipliers_sr_out_r_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_0_Im = multipliers_sr_out_r_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_1_Re = multipliers_sr_out_r_1_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_1_Im = multipliers_sr_out_r_1_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_2_Re = multipliers_sr_out_r_2_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_2_Im = multipliers_sr_out_r_2_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_3_Re = multipliers_sr_out_r_3_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_3_Im = multipliers_sr_out_r_3_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_4_Re = multipliers_sr_out_r_4_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_4_Im = multipliers_sr_out_r_4_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_5_Re = multipliers_sr_out_r_5_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_5_Im = multipliers_sr_out_r_5_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_6_Re = multipliers_sr_out_r_6_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_6_Im = multipliers_sr_out_r_6_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_7_Re = multipliers_sr_out_r_7_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_7_Im = multipliers_sr_out_r_7_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_8_Re = multipliers_sr_out_r_8_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_8_Im = multipliers_sr_out_r_8_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_9_Re = multipliers_sr_out_r_9_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_9_Im = multipliers_sr_out_r_9_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_10_Re = multipliers_sr_out_r_10_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_10_Im = multipliers_sr_out_r_10_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_11_Re = multipliers_sr_out_r_11_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_11_Im = multipliers_sr_out_r_11_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_12_Re = multipliers_sr_out_r_12_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_12_Im = multipliers_sr_out_r_12_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_13_Re = multipliers_sr_out_r_13_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_13_Im = multipliers_sr_out_r_13_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_14_Re = multipliers_sr_out_r_14_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_14_Im = multipliers_sr_out_r_14_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_15_Re = multipliers_sr_out_r_15_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_15_Im = multipliers_sr_out_r_15_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_inv = io_in_inv; // @[TwidFactorDesigns.scala 56:23]
  assign TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_addr = {{4'd0}, value_1}; // @[TwidFactorDesigns.scala 55:24]
  assign FPComplexMultiplier_bw32_clock = clock;
  assign FPComplexMultiplier_bw32_reset = reset;
  assign FPComplexMultiplier_bw32_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_io_in_a_Re = io_in_0_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_io_in_a_Im = io_in_0_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_0_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_1_clock = clock;
  assign FPComplexMultiplier_bw32_1_reset = reset;
  assign FPComplexMultiplier_bw32_1_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_1_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_1_io_in_a_Re = io_in_1_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_1_io_in_a_Im = io_in_1_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_1_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_1_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_1_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_1_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_2_clock = clock;
  assign FPComplexMultiplier_bw32_2_reset = reset;
  assign FPComplexMultiplier_bw32_2_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_2_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_2_io_in_a_Re = io_in_2_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_2_io_in_a_Im = io_in_2_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_2_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_2_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_2_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_3_clock = clock;
  assign FPComplexMultiplier_bw32_3_reset = reset;
  assign FPComplexMultiplier_bw32_3_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_3_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_3_io_in_a_Re = io_in_3_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_3_io_in_a_Im = io_in_3_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_3_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_3_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_3_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_3_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_4_clock = clock;
  assign FPComplexMultiplier_bw32_4_reset = reset;
  assign FPComplexMultiplier_bw32_4_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_4_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_4_io_in_a_Re = io_in_4_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_4_io_in_a_Im = io_in_4_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_4_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_4_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_4_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_5_clock = clock;
  assign FPComplexMultiplier_bw32_5_reset = reset;
  assign FPComplexMultiplier_bw32_5_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_5_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_5_io_in_a_Re = io_in_5_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_5_io_in_a_Im = io_in_5_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_5_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_5_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_5_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_5_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_6_clock = clock;
  assign FPComplexMultiplier_bw32_6_reset = reset;
  assign FPComplexMultiplier_bw32_6_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_6_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_6_io_in_a_Re = io_in_6_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_6_io_in_a_Im = io_in_6_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_6_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_6_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_6_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_7_clock = clock;
  assign FPComplexMultiplier_bw32_7_reset = reset;
  assign FPComplexMultiplier_bw32_7_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_7_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_7_io_in_a_Re = io_in_7_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_7_io_in_a_Im = io_in_7_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_7_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_7_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_7_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_7_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_8_clock = clock;
  assign FPComplexMultiplier_bw32_8_reset = reset;
  assign FPComplexMultiplier_bw32_8_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_8_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_8_io_in_a_Re = io_in_8_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_8_io_in_a_Im = io_in_8_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_8_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_8_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_8_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_9_clock = clock;
  assign FPComplexMultiplier_bw32_9_reset = reset;
  assign FPComplexMultiplier_bw32_9_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_9_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_9_io_in_a_Re = io_in_9_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_9_io_in_a_Im = io_in_9_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_9_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_9_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_9_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_9_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_10_clock = clock;
  assign FPComplexMultiplier_bw32_10_reset = reset;
  assign FPComplexMultiplier_bw32_10_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_10_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_10_io_in_a_Re = io_in_10_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_10_io_in_a_Im = io_in_10_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_10_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_10_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_10_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_11_clock = clock;
  assign FPComplexMultiplier_bw32_11_reset = reset;
  assign FPComplexMultiplier_bw32_11_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_11_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_11_io_in_a_Re = io_in_11_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_11_io_in_a_Im = io_in_11_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_11_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_11_Re
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_11_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_11_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_12_clock = clock;
  assign FPComplexMultiplier_bw32_12_reset = reset;
  assign FPComplexMultiplier_bw32_12_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_12_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_12_io_in_a_Re = io_in_12_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_12_io_in_a_Im = io_in_12_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_12_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_12_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_12_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_13_clock = clock;
  assign FPComplexMultiplier_bw32_13_reset = reset;
  assign FPComplexMultiplier_bw32_13_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_13_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_13_io_in_a_Re = io_in_13_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_13_io_in_a_Im = io_in_13_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_13_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_13_Re
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_13_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_13_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_14_clock = clock;
  assign FPComplexMultiplier_bw32_14_reset = reset;
  assign FPComplexMultiplier_bw32_14_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_14_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_14_io_in_a_Re = io_in_14_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_14_io_in_a_Im = io_in_14_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_14_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_14_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_14_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_15_clock = clock;
  assign FPComplexMultiplier_bw32_15_reset = reset;
  assign FPComplexMultiplier_bw32_15_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_15_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_15_io_in_a_Re = io_in_15_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_15_io_in_a_Im = io_in_15_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_15_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_15_Re
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_15_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_data_15_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en) begin // @[TwidFactorDesigns.scala 57:22]
      if (io_in_valid) begin // @[TwidFactorDesigns.scala 58:27]
        value_1 <= _value_T_1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_Re <= FPComplexMultiplier_bw32_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_Im <= FPComplexMultiplier_bw32_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_1_Re <= FPComplexMultiplier_bw32_1_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_1_Im <= FPComplexMultiplier_bw32_1_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_2_Re <= FPComplexMultiplier_bw32_2_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_2_Im <= FPComplexMultiplier_bw32_2_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_3_Re <= FPComplexMultiplier_bw32_3_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_3_Im <= FPComplexMultiplier_bw32_3_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_4_Re <= FPComplexMultiplier_bw32_4_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_4_Im <= FPComplexMultiplier_bw32_4_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_5_Re <= FPComplexMultiplier_bw32_5_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_5_Im <= FPComplexMultiplier_bw32_5_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_6_Re <= FPComplexMultiplier_bw32_6_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_6_Im <= FPComplexMultiplier_bw32_6_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_7_Re <= FPComplexMultiplier_bw32_7_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_7_Im <= FPComplexMultiplier_bw32_7_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_8_Re <= FPComplexMultiplier_bw32_8_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_8_Im <= FPComplexMultiplier_bw32_8_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_9_Re <= FPComplexMultiplier_bw32_9_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_9_Im <= FPComplexMultiplier_bw32_9_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_10_Re <= FPComplexMultiplier_bw32_10_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_10_Im <= FPComplexMultiplier_bw32_10_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_11_Re <= FPComplexMultiplier_bw32_11_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_11_Im <= FPComplexMultiplier_bw32_11_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_12_Re <= FPComplexMultiplier_bw32_12_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_12_Im <= FPComplexMultiplier_bw32_12_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_13_Re <= FPComplexMultiplier_bw32_13_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_13_Im <= FPComplexMultiplier_bw32_13_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_14_Re <= FPComplexMultiplier_bw32_14_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_14_Im <= FPComplexMultiplier_bw32_14_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_15_Re <= FPComplexMultiplier_bw32_15_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_15_Im <= FPComplexMultiplier_bw32_15_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r <= FPComplexMultiplier_bw32_io_out_valid; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  multipliers_sr_out_r_Re = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  multipliers_sr_out_r_Im = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  multipliers_sr_out_r_1_Re = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  multipliers_sr_out_r_1_Im = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  multipliers_sr_out_r_2_Re = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  multipliers_sr_out_r_2_Im = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  multipliers_sr_out_r_3_Re = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  multipliers_sr_out_r_3_Im = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  multipliers_sr_out_r_4_Re = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  multipliers_sr_out_r_4_Im = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  multipliers_sr_out_r_5_Re = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  multipliers_sr_out_r_5_Im = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  multipliers_sr_out_r_6_Re = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  multipliers_sr_out_r_6_Im = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  multipliers_sr_out_r_7_Re = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  multipliers_sr_out_r_7_Im = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  multipliers_sr_out_r_8_Re = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  multipliers_sr_out_r_8_Im = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  multipliers_sr_out_r_9_Re = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  multipliers_sr_out_r_9_Im = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  multipliers_sr_out_r_10_Re = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  multipliers_sr_out_r_10_Im = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  multipliers_sr_out_r_11_Re = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  multipliers_sr_out_r_11_Im = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  multipliers_sr_out_r_12_Re = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  multipliers_sr_out_r_12_Im = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  multipliers_sr_out_r_13_Re = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  multipliers_sr_out_r_13_Im = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  multipliers_sr_out_r_14_Re = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  multipliers_sr_out_r_14_Im = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  multipliers_sr_out_r_15_Re = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  multipliers_sr_out_r_15_Im = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  io_out_valid_r = _RAND_33[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32(
  input         io_in_inv,
  input  [4:0]  io_in_addr,
  output [31:0] io_out_data_0_Im,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_2_Im,
  output [31:0] io_out_data_3_Re,
  output [31:0] io_out_data_3_Im,
  output [31:0] io_out_data_4_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_6_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im,
  output [31:0] io_out_data_8_Im,
  output [31:0] io_out_data_9_Re,
  output [31:0] io_out_data_9_Im,
  output [31:0] io_out_data_10_Im,
  output [31:0] io_out_data_11_Re,
  output [31:0] io_out_data_11_Im,
  output [31:0] io_out_data_12_Im,
  output [31:0] io_out_data_13_Re,
  output [31:0] io_out_data_13_Im,
  output [31:0] io_out_data_14_Im,
  output [31:0] io_out_data_15_Re,
  output [31:0] io_out_data_15_Im
);
  wire [31:0] _GEN_10 = io_in_addr[0] ? 32'hbe14fdf0 : 32'h3f800000; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_11 = io_in_addr[0] ? 32'h3f7d4694 : 32'h0; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_14 = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_15 = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_26 = io_in_addr[0] ? 32'hbf693fd4 : 32'h3f0a5140; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_27 = io_in_addr[0] ? 32'h3ed30130 : 32'h3f576aa4; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_30 = io_in_addr[0] ? 32'hbe47c5c0 : 32'h3f7b14be; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_31 = io_in_addr[0] ? 32'hbf7b14be : 32'hbe47c5c0; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_42 = io_in_addr[0] ? 32'hbf56cd64 : 32'hbed51130; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_43 = io_in_addr[0] ? 32'hbf0b44f6 : 32'h3f68c7b6; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_46 = io_in_addr[0] ? 32'hbec3ef14 : 32'h3f6c835e; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_47 = io_in_addr[0] ? 32'hbf6c835e : 32'hbec3ef14; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_58 = io_in_addr[0] ? 32'h3b910500 : 32'hbf7d7024; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_59 = io_in_addr[0] ? 32'hbf7fff5a : 32'h3e1081c0; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_62 = io_in_addr[0] ? 32'hbf0e39d8 : 32'h3f54db30; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_63 = io_in_addr[0] ? 32'hbf54db30 : 32'hbf0e39d8; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_74 = io_in_addr[0] ? 32'h3f5806d0 : 32'hbf275530; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_75 = io_in_addr[0] ? 32'hbf095cd6 : 32'hbf41bdce; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_78 = io_in_addr[0] ? 32'hbf3504f2 : 32'h3f3504f2; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_90 = io_in_addr[0] ? 32'h3f684e6e : 32'h3e913c28; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_91 = io_in_addr[0] ? 32'h3ed72020 : 32'hbf757c0e; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_94 = io_in_addr[0] ? 32'hbf54db30 : 32'h3f0e39d8; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_95 = io_in_addr[0] ? 32'hbf0e39d8 : 32'hbf54db30; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_106 = io_in_addr[0] ? 32'h3e0c04d0 : 32'h3f75cdb8; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_107 = io_in_addr[0] ? 32'h3f7d9870 : 32'hbe8f0f8c; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_110 = io_in_addr[0] ? 32'hbf6c835e : 32'h3ec3ef14; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_111 = io_in_addr[0] ? 32'hbec3ef14 : 32'hbf6c835e; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_122 = io_in_addr[0] ? 32'hbf427ae8 : 32'h3f40ffbc; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_123 = io_in_addr[0] ? 32'h3f267942 : 32'h3f283046; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_126 = io_in_addr[0] ? 32'hbf7b14be : 32'h3e47c5c0; // @[TwidFactorDesigns.scala 26:{53,53}]
  wire [31:0] _GEN_127 = io_in_addr[0] ? 32'hbe47c5c0 : 32'hbf7b14be; // @[TwidFactorDesigns.scala 26:{53,53}]
  assign io_out_data_0_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_1_Re = io_in_inv ? _GEN_10 : _GEN_14; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_1_Im = io_in_inv ? _GEN_11 : _GEN_15; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_2_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_3_Re = io_in_inv ? _GEN_26 : _GEN_30; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_3_Im = io_in_inv ? _GEN_27 : _GEN_31; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_4_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_5_Re = io_in_inv ? _GEN_42 : _GEN_46; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_5_Im = io_in_inv ? _GEN_43 : _GEN_47; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_6_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_7_Re = io_in_inv ? _GEN_58 : _GEN_62; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_7_Im = io_in_inv ? _GEN_59 : _GEN_63; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_8_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_9_Re = io_in_inv ? _GEN_74 : _GEN_78; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_9_Im = io_in_inv ? _GEN_75 : 32'hbf3504f2; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_10_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_11_Re = io_in_inv ? _GEN_90 : _GEN_94; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_11_Im = io_in_inv ? _GEN_91 : _GEN_95; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_12_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_13_Re = io_in_inv ? _GEN_106 : _GEN_110; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_13_Im = io_in_inv ? _GEN_107 : _GEN_111; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_14_Im = io_in_inv ? 32'h0 : 32'h80800000; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_15_Re = io_in_inv ? _GEN_122 : _GEN_126; // @[TwidFactorDesigns.scala 26:53]
  assign io_out_data_15_Im = io_in_inv ? _GEN_123 : _GEN_127; // @[TwidFactorDesigns.scala 26:53]
endmodule
module TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32(
  input         clock,
  input         reset,
  input         io_in_inv,
  input         io_in_en,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_valid,
  output        io_out_valid,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  wire  TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_inv; // @[TwidFactorDesigns.scala 49:28]
  wire [4:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_addr; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_0_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_1_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_1_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_2_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_3_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_3_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_4_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_5_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_5_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_6_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_7_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_7_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_8_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_9_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_9_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_10_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_11_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_11_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_12_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_13_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_13_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_14_Im; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_15_Re; // @[TwidFactorDesigns.scala 49:28]
  wire [31:0] TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_15_Im; // @[TwidFactorDesigns.scala 49:28]
  wire  FPComplexMultiplier_bw32_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_1_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_1_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_2_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_2_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_3_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_3_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_4_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_4_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_5_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_5_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_6_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_6_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_7_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_7_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_8_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_8_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_9_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_9_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_10_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_10_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_11_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_11_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_12_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_12_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_13_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_13_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_14_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_14_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_clock; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_reset; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_io_in_en; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_io_in_valid; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_in_a_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_in_a_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_in_b_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_in_b_Im; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_out_s_Re; // @[TwidFactorDesigns.scala 66:48]
  wire [31:0] FPComplexMultiplier_bw32_15_io_out_s_Im; // @[TwidFactorDesigns.scala 66:48]
  wire  FPComplexMultiplier_bw32_15_io_out_valid; // @[TwidFactorDesigns.scala 66:48]
  reg  value_1; // @[Counter.scala 62:40]
  wire  _value_T_1 = value_1 + 1'h1; // @[Counter.scala 78:24]
  reg [31:0] multipliers_sr_out_r_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_1_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_1_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_2_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_2_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_3_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_3_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_4_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_4_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_5_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_5_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_6_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_6_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_7_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_7_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_8_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_8_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_9_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_9_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_10_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_10_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_11_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_11_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_12_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_12_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_13_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_13_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_14_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_14_Im; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_15_Re; // @[Reg.scala 16:16]
  reg [31:0] multipliers_sr_out_r_15_Im; // @[Reg.scala 16:16]
  reg  io_out_valid_r; // @[Reg.scala 16:16]
  TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32 TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32 ( // @[TwidFactorDesigns.scala 49:28]
    .io_in_inv(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_inv),
    .io_in_addr(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_addr),
    .io_out_data_0_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_0_Im),
    .io_out_data_1_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_1_Im),
    .io_out_data_2_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_2_Im),
    .io_out_data_3_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_3_Re),
    .io_out_data_3_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_3_Im),
    .io_out_data_4_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_4_Im),
    .io_out_data_5_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_5_Im),
    .io_out_data_6_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_6_Im),
    .io_out_data_7_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_7_Im),
    .io_out_data_8_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_8_Im),
    .io_out_data_9_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_9_Re),
    .io_out_data_9_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_9_Im),
    .io_out_data_10_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_10_Im),
    .io_out_data_11_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_11_Re),
    .io_out_data_11_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_11_Im),
    .io_out_data_12_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_12_Im),
    .io_out_data_13_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_13_Re),
    .io_out_data_13_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_13_Im),
    .io_out_data_14_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_14_Im),
    .io_out_data_15_Re(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_15_Re),
    .io_out_data_15_Im(TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_15_Im)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_clock),
    .reset(FPComplexMultiplier_bw32_reset),
    .io_in_en(FPComplexMultiplier_bw32_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_1 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_1_clock),
    .reset(FPComplexMultiplier_bw32_1_reset),
    .io_in_en(FPComplexMultiplier_bw32_1_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_1_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_1_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_1_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_2 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_2_clock),
    .reset(FPComplexMultiplier_bw32_2_reset),
    .io_in_en(FPComplexMultiplier_bw32_2_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_2_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_2_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_2_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_3 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_3_clock),
    .reset(FPComplexMultiplier_bw32_3_reset),
    .io_in_en(FPComplexMultiplier_bw32_3_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_3_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_3_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_3_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_4 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_4_clock),
    .reset(FPComplexMultiplier_bw32_4_reset),
    .io_in_en(FPComplexMultiplier_bw32_4_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_4_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_4_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_4_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_5 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_5_clock),
    .reset(FPComplexMultiplier_bw32_5_reset),
    .io_in_en(FPComplexMultiplier_bw32_5_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_5_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_5_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_5_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_6 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_6_clock),
    .reset(FPComplexMultiplier_bw32_6_reset),
    .io_in_en(FPComplexMultiplier_bw32_6_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_6_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_6_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_6_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_7 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_7_clock),
    .reset(FPComplexMultiplier_bw32_7_reset),
    .io_in_en(FPComplexMultiplier_bw32_7_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_7_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_7_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_7_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_8 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_8_clock),
    .reset(FPComplexMultiplier_bw32_8_reset),
    .io_in_en(FPComplexMultiplier_bw32_8_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_8_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_8_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_8_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_8_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_8_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_8_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_9 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_9_clock),
    .reset(FPComplexMultiplier_bw32_9_reset),
    .io_in_en(FPComplexMultiplier_bw32_9_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_9_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_9_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_9_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_10 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_10_clock),
    .reset(FPComplexMultiplier_bw32_10_reset),
    .io_in_en(FPComplexMultiplier_bw32_10_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_10_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_10_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_10_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_10_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_10_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_10_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_11 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_11_clock),
    .reset(FPComplexMultiplier_bw32_11_reset),
    .io_in_en(FPComplexMultiplier_bw32_11_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_11_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_11_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_11_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_12 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_12_clock),
    .reset(FPComplexMultiplier_bw32_12_reset),
    .io_in_en(FPComplexMultiplier_bw32_12_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_12_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_12_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_12_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_12_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_12_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_12_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_13 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_13_clock),
    .reset(FPComplexMultiplier_bw32_13_reset),
    .io_in_en(FPComplexMultiplier_bw32_13_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_13_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_13_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_13_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_14 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_14_clock),
    .reset(FPComplexMultiplier_bw32_14_reset),
    .io_in_en(FPComplexMultiplier_bw32_14_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_14_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_14_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_14_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_14_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_14_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_14_io_out_valid)
  );
  FPComplexMultiplier_bw32 FPComplexMultiplier_bw32_15 ( // @[TwidFactorDesigns.scala 66:48]
    .clock(FPComplexMultiplier_bw32_15_clock),
    .reset(FPComplexMultiplier_bw32_15_reset),
    .io_in_en(FPComplexMultiplier_bw32_15_io_in_en),
    .io_in_valid(FPComplexMultiplier_bw32_15_io_in_valid),
    .io_in_a_Re(FPComplexMultiplier_bw32_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMultiplier_bw32_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMultiplier_bw32_15_io_in_b_Re),
    .io_in_b_Im(FPComplexMultiplier_bw32_15_io_in_b_Im),
    .io_out_s_Re(FPComplexMultiplier_bw32_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMultiplier_bw32_15_io_out_s_Im),
    .io_out_valid(FPComplexMultiplier_bw32_15_io_out_valid)
  );
  assign io_out_valid = io_out_valid_r; // @[TwidFactorDesigns.scala 77:22]
  assign io_out_0_Re = multipliers_sr_out_r_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_0_Im = multipliers_sr_out_r_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_1_Re = multipliers_sr_out_r_1_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_1_Im = multipliers_sr_out_r_1_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_2_Re = multipliers_sr_out_r_2_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_2_Im = multipliers_sr_out_r_2_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_3_Re = multipliers_sr_out_r_3_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_3_Im = multipliers_sr_out_r_3_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_4_Re = multipliers_sr_out_r_4_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_4_Im = multipliers_sr_out_r_4_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_5_Re = multipliers_sr_out_r_5_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_5_Im = multipliers_sr_out_r_5_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_6_Re = multipliers_sr_out_r_6_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_6_Im = multipliers_sr_out_r_6_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_7_Re = multipliers_sr_out_r_7_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_7_Im = multipliers_sr_out_r_7_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_8_Re = multipliers_sr_out_r_8_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_8_Im = multipliers_sr_out_r_8_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_9_Re = multipliers_sr_out_r_9_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_9_Im = multipliers_sr_out_r_9_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_10_Re = multipliers_sr_out_r_10_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_10_Im = multipliers_sr_out_r_10_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_11_Re = multipliers_sr_out_r_11_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_11_Im = multipliers_sr_out_r_11_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_12_Re = multipliers_sr_out_r_12_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_12_Im = multipliers_sr_out_r_12_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_13_Re = multipliers_sr_out_r_13_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_13_Im = multipliers_sr_out_r_13_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_14_Re = multipliers_sr_out_r_14_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_14_Im = multipliers_sr_out_r_14_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_15_Re = multipliers_sr_out_r_15_Re; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign io_out_15_Im = multipliers_sr_out_r_15_Im; // @[TwidFactorDesigns.scala 73:{41,41}]
  assign TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_inv = io_in_inv; // @[TwidFactorDesigns.scala 56:23]
  assign TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_addr = {{4'd0}, value_1}; // @[TwidFactorDesigns.scala 55:24]
  assign FPComplexMultiplier_bw32_clock = clock;
  assign FPComplexMultiplier_bw32_reset = reset;
  assign FPComplexMultiplier_bw32_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_io_in_a_Re = io_in_0_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_io_in_a_Im = io_in_0_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_0_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_1_clock = clock;
  assign FPComplexMultiplier_bw32_1_reset = reset;
  assign FPComplexMultiplier_bw32_1_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_1_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_1_io_in_a_Re = io_in_1_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_1_io_in_a_Im = io_in_1_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_1_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_1_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_1_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_1_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_2_clock = clock;
  assign FPComplexMultiplier_bw32_2_reset = reset;
  assign FPComplexMultiplier_bw32_2_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_2_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_2_io_in_a_Re = io_in_2_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_2_io_in_a_Im = io_in_2_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_2_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_2_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_2_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_3_clock = clock;
  assign FPComplexMultiplier_bw32_3_reset = reset;
  assign FPComplexMultiplier_bw32_3_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_3_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_3_io_in_a_Re = io_in_3_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_3_io_in_a_Im = io_in_3_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_3_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_3_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_3_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_3_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_4_clock = clock;
  assign FPComplexMultiplier_bw32_4_reset = reset;
  assign FPComplexMultiplier_bw32_4_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_4_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_4_io_in_a_Re = io_in_4_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_4_io_in_a_Im = io_in_4_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_4_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_4_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_4_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_5_clock = clock;
  assign FPComplexMultiplier_bw32_5_reset = reset;
  assign FPComplexMultiplier_bw32_5_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_5_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_5_io_in_a_Re = io_in_5_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_5_io_in_a_Im = io_in_5_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_5_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_5_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_5_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_5_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_6_clock = clock;
  assign FPComplexMultiplier_bw32_6_reset = reset;
  assign FPComplexMultiplier_bw32_6_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_6_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_6_io_in_a_Re = io_in_6_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_6_io_in_a_Im = io_in_6_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_6_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_6_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_6_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_7_clock = clock;
  assign FPComplexMultiplier_bw32_7_reset = reset;
  assign FPComplexMultiplier_bw32_7_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_7_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_7_io_in_a_Re = io_in_7_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_7_io_in_a_Im = io_in_7_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_7_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_7_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_7_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_7_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_8_clock = clock;
  assign FPComplexMultiplier_bw32_8_reset = reset;
  assign FPComplexMultiplier_bw32_8_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_8_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_8_io_in_a_Re = io_in_8_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_8_io_in_a_Im = io_in_8_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_8_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_8_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_8_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_9_clock = clock;
  assign FPComplexMultiplier_bw32_9_reset = reset;
  assign FPComplexMultiplier_bw32_9_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_9_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_9_io_in_a_Re = io_in_9_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_9_io_in_a_Im = io_in_9_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_9_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_9_Re; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_9_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_9_Im; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_10_clock = clock;
  assign FPComplexMultiplier_bw32_10_reset = reset;
  assign FPComplexMultiplier_bw32_10_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_10_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_10_io_in_a_Re = io_in_10_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_10_io_in_a_Im = io_in_10_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_10_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_10_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_10_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_11_clock = clock;
  assign FPComplexMultiplier_bw32_11_reset = reset;
  assign FPComplexMultiplier_bw32_11_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_11_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_11_io_in_a_Re = io_in_11_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_11_io_in_a_Im = io_in_11_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_11_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_11_Re
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_11_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_11_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_12_clock = clock;
  assign FPComplexMultiplier_bw32_12_reset = reset;
  assign FPComplexMultiplier_bw32_12_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_12_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_12_io_in_a_Re = io_in_12_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_12_io_in_a_Im = io_in_12_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_12_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_12_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_12_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_13_clock = clock;
  assign FPComplexMultiplier_bw32_13_reset = reset;
  assign FPComplexMultiplier_bw32_13_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_13_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_13_io_in_a_Re = io_in_13_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_13_io_in_a_Im = io_in_13_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_13_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_13_Re
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_13_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_13_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_14_clock = clock;
  assign FPComplexMultiplier_bw32_14_reset = reset;
  assign FPComplexMultiplier_bw32_14_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_14_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_14_io_in_a_Re = io_in_14_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_14_io_in_a_Im = io_in_14_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_14_io_in_b_Re = 32'h3f800000; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_14_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_14_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_15_clock = clock;
  assign FPComplexMultiplier_bw32_15_reset = reset;
  assign FPComplexMultiplier_bw32_15_io_in_en = io_in_en; // @[TwidFactorDesigns.scala 69:32]
  assign FPComplexMultiplier_bw32_15_io_in_valid = io_in_valid; // @[TwidFactorDesigns.scala 68:35]
  assign FPComplexMultiplier_bw32_15_io_in_a_Re = io_in_15_Re; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_15_io_in_a_Im = io_in_15_Im; // @[TwidFactorDesigns.scala 70:31]
  assign FPComplexMultiplier_bw32_15_io_in_b_Re = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_15_Re
    ; // @[TwidFactorDesigns.scala 71:31]
  assign FPComplexMultiplier_bw32_15_io_in_b_Im = TwiddleFactorROM_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_data_15_Im
    ; // @[TwidFactorDesigns.scala 71:31]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_in_en) begin // @[TwidFactorDesigns.scala 57:22]
      if (io_in_valid) begin // @[TwidFactorDesigns.scala 58:27]
        value_1 <= _value_T_1;
      end
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_Re <= FPComplexMultiplier_bw32_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_Im <= FPComplexMultiplier_bw32_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_1_Re <= FPComplexMultiplier_bw32_1_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_1_Im <= FPComplexMultiplier_bw32_1_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_2_Re <= FPComplexMultiplier_bw32_2_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_2_Im <= FPComplexMultiplier_bw32_2_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_3_Re <= FPComplexMultiplier_bw32_3_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_3_Im <= FPComplexMultiplier_bw32_3_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_4_Re <= FPComplexMultiplier_bw32_4_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_4_Im <= FPComplexMultiplier_bw32_4_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_5_Re <= FPComplexMultiplier_bw32_5_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_5_Im <= FPComplexMultiplier_bw32_5_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_6_Re <= FPComplexMultiplier_bw32_6_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_6_Im <= FPComplexMultiplier_bw32_6_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_7_Re <= FPComplexMultiplier_bw32_7_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_7_Im <= FPComplexMultiplier_bw32_7_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_8_Re <= FPComplexMultiplier_bw32_8_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_8_Im <= FPComplexMultiplier_bw32_8_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_9_Re <= FPComplexMultiplier_bw32_9_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_9_Im <= FPComplexMultiplier_bw32_9_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_10_Re <= FPComplexMultiplier_bw32_10_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_10_Im <= FPComplexMultiplier_bw32_10_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_11_Re <= FPComplexMultiplier_bw32_11_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_11_Im <= FPComplexMultiplier_bw32_11_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_12_Re <= FPComplexMultiplier_bw32_12_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_12_Im <= FPComplexMultiplier_bw32_12_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_13_Re <= FPComplexMultiplier_bw32_13_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_13_Im <= FPComplexMultiplier_bw32_13_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_14_Re <= FPComplexMultiplier_bw32_14_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_14_Im <= FPComplexMultiplier_bw32_14_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_15_Re <= FPComplexMultiplier_bw32_15_io_out_s_Re; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      multipliers_sr_out_r_15_Im <= FPComplexMultiplier_bw32_15_io_out_s_Im; // @[Reg.scala 17:22]
    end
    if (io_in_en) begin // @[Reg.scala 17:18]
      io_out_valid_r <= FPComplexMultiplier_bw32_io_out_valid; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  multipliers_sr_out_r_Re = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  multipliers_sr_out_r_Im = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  multipliers_sr_out_r_1_Re = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  multipliers_sr_out_r_1_Im = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  multipliers_sr_out_r_2_Re = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  multipliers_sr_out_r_2_Im = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  multipliers_sr_out_r_3_Re = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  multipliers_sr_out_r_3_Im = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  multipliers_sr_out_r_4_Re = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  multipliers_sr_out_r_4_Im = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  multipliers_sr_out_r_5_Re = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  multipliers_sr_out_r_5_Im = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  multipliers_sr_out_r_6_Re = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  multipliers_sr_out_r_6_Im = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  multipliers_sr_out_r_7_Re = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  multipliers_sr_out_r_7_Im = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  multipliers_sr_out_r_8_Re = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  multipliers_sr_out_r_8_Im = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  multipliers_sr_out_r_9_Re = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  multipliers_sr_out_r_9_Im = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  multipliers_sr_out_r_10_Re = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  multipliers_sr_out_r_10_Im = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  multipliers_sr_out_r_11_Re = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  multipliers_sr_out_r_11_Im = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  multipliers_sr_out_r_12_Re = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  multipliers_sr_out_r_12_Im = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  multipliers_sr_out_r_13_Re = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  multipliers_sr_out_r_13_Im = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  multipliers_sr_out_r_14_Re = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  multipliers_sr_out_r_14_Im = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  multipliers_sr_out_r_15_Re = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  multipliers_sr_out_r_15_Im = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  io_out_valid_r = _RAND_33[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FFT32w16(
  input         clock,
  input         reset,
  input         io_in_inv,
  input         io_in_ready,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_valid,
  output        io_out_valid,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output        io_out_ready
);
  wire  DFT2_bw32_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_1_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_1_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_1_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_1_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_1_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_1_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_1_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_1_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_1_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_1_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_1_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_1_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_1_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_2_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_2_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_2_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_2_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_2_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_2_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_2_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_2_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_2_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_2_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_2_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_2_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_2_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_3_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_3_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_3_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_3_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_3_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_3_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_3_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_3_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_3_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_3_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_3_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_3_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_3_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_4_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_4_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_4_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_4_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_4_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_4_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_4_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_4_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_4_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_4_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_4_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_4_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_4_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_5_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_5_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_5_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_5_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_5_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_5_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_5_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_5_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_5_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_5_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_5_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_5_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_5_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_6_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_6_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_6_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_6_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_6_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_6_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_6_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_6_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_6_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_6_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_6_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_6_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_6_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_7_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_7_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_7_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_7_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_7_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_7_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_7_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_7_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_7_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_7_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_7_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_7_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_7_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_8_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_8_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_8_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_8_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_8_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_8_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_8_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_8_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_8_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_8_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_8_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_8_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_8_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_9_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_9_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_9_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_9_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_9_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_9_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_9_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_9_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_9_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_9_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_9_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_9_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_9_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_10_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_10_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_10_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_10_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_10_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_10_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_10_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_10_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_10_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_10_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_10_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_10_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_10_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_11_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_11_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_11_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_11_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_11_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_11_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_11_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_11_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_11_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_11_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_11_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_11_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_11_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_12_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_12_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_12_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_12_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_12_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_12_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_12_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_12_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_12_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_12_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_12_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_12_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_12_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_13_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_13_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_13_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_13_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_13_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_13_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_13_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_13_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_13_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_13_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_13_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_13_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_13_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_14_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_14_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_14_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_14_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_14_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_14_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_14_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_14_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_14_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_14_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_14_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_14_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_14_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_15_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_15_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_15_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_15_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_15_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_15_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_15_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_15_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_15_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_15_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_15_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_15_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_15_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_16_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_16_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_16_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_16_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_16_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_16_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_16_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_16_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_16_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_16_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_16_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_16_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_16_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_17_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_17_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_17_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_17_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_17_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_17_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_17_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_17_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_17_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_17_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_17_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_17_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_17_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_18_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_18_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_18_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_18_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_18_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_18_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_18_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_18_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_18_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_18_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_18_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_18_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_18_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_19_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_19_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_19_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_19_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_19_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_19_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_19_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_19_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_19_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_19_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_19_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_19_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_19_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_20_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_20_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_20_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_20_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_20_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_20_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_20_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_20_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_20_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_20_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_20_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_20_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_20_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_21_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_21_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_21_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_21_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_21_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_21_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_21_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_21_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_21_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_21_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_21_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_21_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_21_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_22_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_22_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_22_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_22_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_22_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_22_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_22_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_22_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_22_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_22_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_22_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_22_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_22_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_23_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_23_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_23_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_23_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_23_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_23_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_23_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_23_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_23_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_23_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_23_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_23_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_23_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_24_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_24_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_24_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_24_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_24_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_24_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_24_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_24_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_24_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_24_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_24_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_24_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_24_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_25_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_25_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_25_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_25_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_25_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_25_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_25_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_25_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_25_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_25_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_25_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_25_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_25_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_26_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_26_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_26_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_26_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_26_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_26_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_26_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_26_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_26_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_26_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_26_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_26_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_26_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_27_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_27_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_27_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_27_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_27_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_27_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_27_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_27_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_27_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_27_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_27_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_27_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_27_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_28_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_28_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_28_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_28_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_28_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_28_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_28_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_28_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_28_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_28_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_28_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_28_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_28_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_29_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_29_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_29_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_29_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_29_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_29_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_29_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_29_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_29_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_29_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_29_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_29_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_29_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_30_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_30_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_30_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_30_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_30_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_30_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_30_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_30_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_30_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_30_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_30_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_30_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_30_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_31_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_31_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_31_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_31_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_31_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_31_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_31_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_31_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_31_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_31_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_31_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_31_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_31_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_32_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_32_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_32_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_32_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_32_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_32_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_32_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_32_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_32_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_32_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_32_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_32_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_32_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_33_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_33_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_33_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_33_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_33_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_33_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_33_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_33_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_33_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_33_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_33_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_33_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_33_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_34_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_34_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_34_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_34_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_34_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_34_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_34_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_34_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_34_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_34_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_34_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_34_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_34_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_35_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_35_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_35_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_35_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_35_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_35_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_35_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_35_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_35_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_35_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_35_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_35_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_35_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_36_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_36_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_36_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_36_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_36_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_36_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_36_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_36_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_36_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_36_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_36_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_36_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_36_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_37_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_37_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_37_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_37_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_37_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_37_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_37_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_37_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_37_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_37_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_37_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_37_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_37_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_38_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_38_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_38_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_38_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_38_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_38_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_38_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_38_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_38_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_38_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_38_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_38_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_38_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_39_clock; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_39_reset; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_39_io_in_en; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_39_io_in_valid; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_39_io_in_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_39_io_in_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_39_io_in_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_39_io_in_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_39_io_out_0_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_39_io_out_0_Im; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_39_io_out_1_Re; // @[FFTSRDesigns.scala 79:70]
  wire [31:0] DFT2_bw32_39_io_out_1_Im; // @[FFTSRDesigns.scala 79:70]
  wire  DFT2_bw32_39_io_out_valid; // @[FFTSRDesigns.scala 79:70]
  wire  Permute_Streaming_N32_r2_w16_bitRtrue_bw64_clock; // @[FFTSRDesigns.scala 82:15]
  wire  Permute_Streaming_N32_r2_w16_bitRtrue_bw64_reset; // @[FFTSRDesigns.scala 82:15]
  wire  Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_en; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_0; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_1; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_2; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_3; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_4; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_5; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_6; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_7; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_8; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_9; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_10; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_11; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_12; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_13; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_14; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_15; // @[FFTSRDesigns.scala 82:15]
  wire  Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_valid; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_0; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_1; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_2; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_3; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_4; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_5; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_6; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_7; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_8; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_9; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_10; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_11; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_12; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_13; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_14; // @[FFTSRDesigns.scala 82:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_15; // @[FFTSRDesigns.scala 82:15]
  wire  Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_valid; // @[FFTSRDesigns.scala 82:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_clock; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_reset; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_en; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_0; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_1; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_2; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_3; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_4; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_5; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_6; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_7; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_8; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_9; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_10; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_11; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_12; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_13; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_14; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_15; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_valid; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_0; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_1; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_2; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_3; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_4; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_5; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_6; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_7; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_8; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_9; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_10; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_11; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_12; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_13; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_14; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_15; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_valid; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_clock; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_reset; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_en; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_0; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_1; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_2; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_3; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_4; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_5; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_6; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_7; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_8; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_9; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_10; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_11; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_12; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_13; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_14; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_15; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_valid; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_0; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_1; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_2; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_3; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_4; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_5; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_6; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_7; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_8; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_9; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_10; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_11; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_12; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_13; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_14; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_15; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_valid; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_clock; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_reset; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_en; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_0; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_1; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_2; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_3; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_4; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_5; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_6; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_7; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_8; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_9; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_10; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_11; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_12; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_13; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_14; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_15; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_valid; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_0; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_1; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_2; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_3; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_4; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_5; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_6; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_7; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_8; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_9; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_10; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_11; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_12; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_13; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_14; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_15; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_valid; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_clock; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_reset; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_en; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_0; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_1; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_2; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_3; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_4; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_5; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_6; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_7; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_8; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_9; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_10; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_11; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_12; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_13; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_14; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_15; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_valid; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_0; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_1; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_2; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_3; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_4; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_5; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_6; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_7; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_8; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_9; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_10; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_11; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_12; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_13; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_14; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_15; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_valid; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_clock; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_reset; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_en; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_0; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_1; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_2; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_3; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_4; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_5; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_6; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_7; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_8; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_9; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_10; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_11; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_12; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_13; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_14; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_15; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_valid; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_0; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_1; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_2; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_3; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_4; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_5; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_6; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_7; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_8; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_9; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_10; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_11; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_12; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_13; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_14; // @[FFTSRDesigns.scala 84:15]
  wire [63:0] Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_15; // @[FFTSRDesigns.scala 84:15]
  wire  Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_valid; // @[FFTSRDesigns.scala 84:15]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_clock; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_reset; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_inv; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_en; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_0_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_0_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_1_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_1_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_2_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_2_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_3_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_3_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_4_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_4_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_5_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_5_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_6_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_6_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_7_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_7_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_8_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_8_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_9_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_9_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_10_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_10_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_11_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_11_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_12_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_12_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_13_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_13_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_14_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_14_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_15_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_15_Im; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_valid; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_valid; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_0_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_0_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_1_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_1_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_2_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_2_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_3_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_3_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_4_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_4_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_5_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_5_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_6_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_6_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_7_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_7_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_8_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_8_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_9_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_9_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_10_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_10_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_11_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_11_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_12_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_12_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_13_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_13_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_14_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_14_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_15_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_15_Im; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_clock; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_reset; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_inv; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_en; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_0_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_0_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_1_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_1_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_2_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_2_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_3_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_3_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_4_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_4_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_5_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_5_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_6_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_6_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_7_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_7_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_8_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_8_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_9_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_9_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_10_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_10_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_11_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_11_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_12_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_12_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_13_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_13_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_14_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_14_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_15_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_15_Im; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_valid; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_valid; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_0_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_0_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_1_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_1_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_2_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_2_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_3_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_3_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_4_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_4_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_5_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_5_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_6_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_6_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_7_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_7_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_8_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_8_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_9_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_9_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_10_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_10_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_11_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_11_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_12_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_12_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_13_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_13_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_14_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_14_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_15_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_15_Im; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_clock; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_reset; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_inv; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_en; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_0_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_0_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_1_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_1_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_2_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_2_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_3_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_3_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_4_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_4_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_5_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_5_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_6_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_6_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_7_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_7_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_8_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_8_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_9_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_9_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_10_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_10_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_11_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_11_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_12_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_12_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_13_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_13_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_14_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_14_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_15_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_15_Im; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_valid; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_valid; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_0_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_0_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_1_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_1_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_2_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_2_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_3_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_3_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_4_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_4_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_5_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_5_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_6_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_6_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_7_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_7_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_8_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_8_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_9_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_9_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_10_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_10_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_11_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_11_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_12_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_12_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_13_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_13_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_14_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_14_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_15_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_15_Im; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_clock; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_reset; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_inv; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_en; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_0_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_0_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_1_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_1_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_2_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_2_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_3_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_3_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_4_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_4_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_5_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_5_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_6_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_6_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_7_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_7_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_8_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_8_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_9_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_9_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_10_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_10_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_11_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_11_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_12_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_12_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_13_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_13_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_14_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_14_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_15_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_15_Im; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_valid; // @[FFTSRDesigns.scala 86:68]
  wire  TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_valid; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_0_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_0_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_1_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_1_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_2_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_2_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_3_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_3_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_4_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_4_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_5_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_5_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_6_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_6_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_7_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_7_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_8_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_8_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_9_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_9_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_10_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_10_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_11_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_11_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_12_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_12_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_13_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_13_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_14_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_14_Im; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_15_Re; // @[FFTSRDesigns.scala 86:68]
  wire [31:0] TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_15_Im; // @[FFTSRDesigns.scala 86:68]
  wire [63:0] _WIRE_1 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_0;
  wire [63:0] _WIRE_3 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_1;
  wire [63:0] _WIRE_5 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_2;
  wire [63:0] _WIRE_7 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_3;
  wire [63:0] _WIRE_9 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_4;
  wire [63:0] _WIRE_11 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_5;
  wire [63:0] _WIRE_13 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_6;
  wire [63:0] _WIRE_15 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_7;
  wire [63:0] _WIRE_17 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_8;
  wire [63:0] _WIRE_19 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_9;
  wire [63:0] _WIRE_21 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_10;
  wire [63:0] _WIRE_23 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_11;
  wire [63:0] _WIRE_25 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_12;
  wire [63:0] _WIRE_27 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_13;
  wire [63:0] _WIRE_29 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_14;
  wire [63:0] _WIRE_31 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_15;
  wire [63:0] _WIRE_44 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_0;
  wire [63:0] _WIRE_46 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_1;
  wire [63:0] _WIRE_49 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_2;
  wire [63:0] _WIRE_51 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_3;
  wire [63:0] _WIRE_54 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_4;
  wire [63:0] _WIRE_56 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_5;
  wire [63:0] _WIRE_59 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_6;
  wire [63:0] _WIRE_61 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_7;
  wire [63:0] _WIRE_64 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_8;
  wire [63:0] _WIRE_66 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_9;
  wire [63:0] _WIRE_69 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_10;
  wire [63:0] _WIRE_71 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_11;
  wire [63:0] _WIRE_74 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_12;
  wire [63:0] _WIRE_76 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_13;
  wire [63:0] _WIRE_79 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_14;
  wire [63:0] _WIRE_81 = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_15;
  wire [63:0] _WIRE_93 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_0;
  wire [63:0] _WIRE_95 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_1;
  wire [63:0] _WIRE_97 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_2;
  wire [63:0] _WIRE_99 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_3;
  wire [63:0] _WIRE_101 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_4;
  wire [63:0] _WIRE_103 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_5;
  wire [63:0] _WIRE_105 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_6;
  wire [63:0] _WIRE_107 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_7;
  wire [63:0] _WIRE_109 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_8;
  wire [63:0] _WIRE_111 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_9;
  wire [63:0] _WIRE_113 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_10;
  wire [63:0] _WIRE_115 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_11;
  wire [63:0] _WIRE_117 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_12;
  wire [63:0] _WIRE_119 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_13;
  wire [63:0] _WIRE_121 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_14;
  wire [63:0] _WIRE_123 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_15;
  wire [63:0] _WIRE_143 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_0;
  wire [63:0] _WIRE_145 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_1;
  wire [63:0] _WIRE_147 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_2;
  wire [63:0] _WIRE_149 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_3;
  wire [63:0] _WIRE_151 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_4;
  wire [63:0] _WIRE_153 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_5;
  wire [63:0] _WIRE_155 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_6;
  wire [63:0] _WIRE_157 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_7;
  wire [63:0] _WIRE_159 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_8;
  wire [63:0] _WIRE_161 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_9;
  wire [63:0] _WIRE_163 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_10;
  wire [63:0] _WIRE_165 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_11;
  wire [63:0] _WIRE_167 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_12;
  wire [63:0] _WIRE_169 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_13;
  wire [63:0] _WIRE_171 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_14;
  wire [63:0] _WIRE_173 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_15;
  wire [63:0] _WIRE_193 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_0;
  wire [63:0] _WIRE_195 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_1;
  wire [63:0] _WIRE_197 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_2;
  wire [63:0] _WIRE_199 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_3;
  wire [63:0] _WIRE_201 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_4;
  wire [63:0] _WIRE_203 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_5;
  wire [63:0] _WIRE_205 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_6;
  wire [63:0] _WIRE_207 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_7;
  wire [63:0] _WIRE_209 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_8;
  wire [63:0] _WIRE_211 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_9;
  wire [63:0] _WIRE_213 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_10;
  wire [63:0] _WIRE_215 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_11;
  wire [63:0] _WIRE_217 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_12;
  wire [63:0] _WIRE_219 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_13;
  wire [63:0] _WIRE_221 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_14;
  wire [63:0] _WIRE_223 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_15;
  wire [63:0] _WIRE_243 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_0;
  wire [63:0] _WIRE_245 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_1;
  wire [63:0] _WIRE_247 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_2;
  wire [63:0] _WIRE_249 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_3;
  wire [63:0] _WIRE_251 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_4;
  wire [63:0] _WIRE_253 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_5;
  wire [63:0] _WIRE_255 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_6;
  wire [63:0] _WIRE_257 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_7;
  wire [63:0] _WIRE_259 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_8;
  wire [63:0] _WIRE_261 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_9;
  wire [63:0] _WIRE_263 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_10;
  wire [63:0] _WIRE_265 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_11;
  wire [63:0] _WIRE_267 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_12;
  wire [63:0] _WIRE_269 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_13;
  wire [63:0] _WIRE_271 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_14;
  wire [63:0] _WIRE_273 = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_15;
  DFT2_bw32 DFT2_bw32 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_clock),
    .reset(DFT2_bw32_reset),
    .io_in_en(DFT2_bw32_io_in_en),
    .io_in_valid(DFT2_bw32_io_in_valid),
    .io_in_0_Re(DFT2_bw32_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_io_out_1_Im),
    .io_out_valid(DFT2_bw32_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_1 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_1_clock),
    .reset(DFT2_bw32_1_reset),
    .io_in_en(DFT2_bw32_1_io_in_en),
    .io_in_valid(DFT2_bw32_1_io_in_valid),
    .io_in_0_Re(DFT2_bw32_1_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_1_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_1_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_1_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_1_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_1_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_1_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_1_io_out_1_Im),
    .io_out_valid(DFT2_bw32_1_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_2 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_2_clock),
    .reset(DFT2_bw32_2_reset),
    .io_in_en(DFT2_bw32_2_io_in_en),
    .io_in_valid(DFT2_bw32_2_io_in_valid),
    .io_in_0_Re(DFT2_bw32_2_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_2_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_2_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_2_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_2_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_2_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_2_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_2_io_out_1_Im),
    .io_out_valid(DFT2_bw32_2_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_3 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_3_clock),
    .reset(DFT2_bw32_3_reset),
    .io_in_en(DFT2_bw32_3_io_in_en),
    .io_in_valid(DFT2_bw32_3_io_in_valid),
    .io_in_0_Re(DFT2_bw32_3_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_3_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_3_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_3_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_3_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_3_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_3_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_3_io_out_1_Im),
    .io_out_valid(DFT2_bw32_3_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_4 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_4_clock),
    .reset(DFT2_bw32_4_reset),
    .io_in_en(DFT2_bw32_4_io_in_en),
    .io_in_valid(DFT2_bw32_4_io_in_valid),
    .io_in_0_Re(DFT2_bw32_4_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_4_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_4_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_4_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_4_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_4_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_4_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_4_io_out_1_Im),
    .io_out_valid(DFT2_bw32_4_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_5 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_5_clock),
    .reset(DFT2_bw32_5_reset),
    .io_in_en(DFT2_bw32_5_io_in_en),
    .io_in_valid(DFT2_bw32_5_io_in_valid),
    .io_in_0_Re(DFT2_bw32_5_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_5_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_5_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_5_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_5_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_5_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_5_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_5_io_out_1_Im),
    .io_out_valid(DFT2_bw32_5_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_6 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_6_clock),
    .reset(DFT2_bw32_6_reset),
    .io_in_en(DFT2_bw32_6_io_in_en),
    .io_in_valid(DFT2_bw32_6_io_in_valid),
    .io_in_0_Re(DFT2_bw32_6_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_6_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_6_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_6_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_6_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_6_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_6_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_6_io_out_1_Im),
    .io_out_valid(DFT2_bw32_6_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_7 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_7_clock),
    .reset(DFT2_bw32_7_reset),
    .io_in_en(DFT2_bw32_7_io_in_en),
    .io_in_valid(DFT2_bw32_7_io_in_valid),
    .io_in_0_Re(DFT2_bw32_7_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_7_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_7_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_7_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_7_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_7_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_7_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_7_io_out_1_Im),
    .io_out_valid(DFT2_bw32_7_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_8 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_8_clock),
    .reset(DFT2_bw32_8_reset),
    .io_in_en(DFT2_bw32_8_io_in_en),
    .io_in_valid(DFT2_bw32_8_io_in_valid),
    .io_in_0_Re(DFT2_bw32_8_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_8_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_8_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_8_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_8_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_8_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_8_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_8_io_out_1_Im),
    .io_out_valid(DFT2_bw32_8_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_9 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_9_clock),
    .reset(DFT2_bw32_9_reset),
    .io_in_en(DFT2_bw32_9_io_in_en),
    .io_in_valid(DFT2_bw32_9_io_in_valid),
    .io_in_0_Re(DFT2_bw32_9_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_9_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_9_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_9_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_9_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_9_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_9_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_9_io_out_1_Im),
    .io_out_valid(DFT2_bw32_9_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_10 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_10_clock),
    .reset(DFT2_bw32_10_reset),
    .io_in_en(DFT2_bw32_10_io_in_en),
    .io_in_valid(DFT2_bw32_10_io_in_valid),
    .io_in_0_Re(DFT2_bw32_10_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_10_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_10_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_10_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_10_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_10_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_10_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_10_io_out_1_Im),
    .io_out_valid(DFT2_bw32_10_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_11 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_11_clock),
    .reset(DFT2_bw32_11_reset),
    .io_in_en(DFT2_bw32_11_io_in_en),
    .io_in_valid(DFT2_bw32_11_io_in_valid),
    .io_in_0_Re(DFT2_bw32_11_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_11_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_11_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_11_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_11_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_11_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_11_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_11_io_out_1_Im),
    .io_out_valid(DFT2_bw32_11_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_12 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_12_clock),
    .reset(DFT2_bw32_12_reset),
    .io_in_en(DFT2_bw32_12_io_in_en),
    .io_in_valid(DFT2_bw32_12_io_in_valid),
    .io_in_0_Re(DFT2_bw32_12_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_12_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_12_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_12_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_12_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_12_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_12_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_12_io_out_1_Im),
    .io_out_valid(DFT2_bw32_12_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_13 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_13_clock),
    .reset(DFT2_bw32_13_reset),
    .io_in_en(DFT2_bw32_13_io_in_en),
    .io_in_valid(DFT2_bw32_13_io_in_valid),
    .io_in_0_Re(DFT2_bw32_13_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_13_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_13_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_13_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_13_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_13_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_13_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_13_io_out_1_Im),
    .io_out_valid(DFT2_bw32_13_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_14 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_14_clock),
    .reset(DFT2_bw32_14_reset),
    .io_in_en(DFT2_bw32_14_io_in_en),
    .io_in_valid(DFT2_bw32_14_io_in_valid),
    .io_in_0_Re(DFT2_bw32_14_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_14_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_14_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_14_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_14_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_14_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_14_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_14_io_out_1_Im),
    .io_out_valid(DFT2_bw32_14_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_15 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_15_clock),
    .reset(DFT2_bw32_15_reset),
    .io_in_en(DFT2_bw32_15_io_in_en),
    .io_in_valid(DFT2_bw32_15_io_in_valid),
    .io_in_0_Re(DFT2_bw32_15_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_15_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_15_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_15_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_15_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_15_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_15_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_15_io_out_1_Im),
    .io_out_valid(DFT2_bw32_15_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_16 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_16_clock),
    .reset(DFT2_bw32_16_reset),
    .io_in_en(DFT2_bw32_16_io_in_en),
    .io_in_valid(DFT2_bw32_16_io_in_valid),
    .io_in_0_Re(DFT2_bw32_16_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_16_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_16_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_16_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_16_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_16_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_16_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_16_io_out_1_Im),
    .io_out_valid(DFT2_bw32_16_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_17 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_17_clock),
    .reset(DFT2_bw32_17_reset),
    .io_in_en(DFT2_bw32_17_io_in_en),
    .io_in_valid(DFT2_bw32_17_io_in_valid),
    .io_in_0_Re(DFT2_bw32_17_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_17_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_17_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_17_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_17_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_17_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_17_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_17_io_out_1_Im),
    .io_out_valid(DFT2_bw32_17_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_18 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_18_clock),
    .reset(DFT2_bw32_18_reset),
    .io_in_en(DFT2_bw32_18_io_in_en),
    .io_in_valid(DFT2_bw32_18_io_in_valid),
    .io_in_0_Re(DFT2_bw32_18_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_18_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_18_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_18_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_18_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_18_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_18_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_18_io_out_1_Im),
    .io_out_valid(DFT2_bw32_18_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_19 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_19_clock),
    .reset(DFT2_bw32_19_reset),
    .io_in_en(DFT2_bw32_19_io_in_en),
    .io_in_valid(DFT2_bw32_19_io_in_valid),
    .io_in_0_Re(DFT2_bw32_19_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_19_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_19_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_19_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_19_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_19_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_19_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_19_io_out_1_Im),
    .io_out_valid(DFT2_bw32_19_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_20 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_20_clock),
    .reset(DFT2_bw32_20_reset),
    .io_in_en(DFT2_bw32_20_io_in_en),
    .io_in_valid(DFT2_bw32_20_io_in_valid),
    .io_in_0_Re(DFT2_bw32_20_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_20_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_20_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_20_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_20_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_20_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_20_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_20_io_out_1_Im),
    .io_out_valid(DFT2_bw32_20_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_21 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_21_clock),
    .reset(DFT2_bw32_21_reset),
    .io_in_en(DFT2_bw32_21_io_in_en),
    .io_in_valid(DFT2_bw32_21_io_in_valid),
    .io_in_0_Re(DFT2_bw32_21_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_21_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_21_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_21_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_21_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_21_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_21_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_21_io_out_1_Im),
    .io_out_valid(DFT2_bw32_21_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_22 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_22_clock),
    .reset(DFT2_bw32_22_reset),
    .io_in_en(DFT2_bw32_22_io_in_en),
    .io_in_valid(DFT2_bw32_22_io_in_valid),
    .io_in_0_Re(DFT2_bw32_22_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_22_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_22_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_22_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_22_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_22_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_22_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_22_io_out_1_Im),
    .io_out_valid(DFT2_bw32_22_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_23 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_23_clock),
    .reset(DFT2_bw32_23_reset),
    .io_in_en(DFT2_bw32_23_io_in_en),
    .io_in_valid(DFT2_bw32_23_io_in_valid),
    .io_in_0_Re(DFT2_bw32_23_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_23_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_23_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_23_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_23_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_23_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_23_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_23_io_out_1_Im),
    .io_out_valid(DFT2_bw32_23_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_24 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_24_clock),
    .reset(DFT2_bw32_24_reset),
    .io_in_en(DFT2_bw32_24_io_in_en),
    .io_in_valid(DFT2_bw32_24_io_in_valid),
    .io_in_0_Re(DFT2_bw32_24_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_24_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_24_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_24_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_24_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_24_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_24_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_24_io_out_1_Im),
    .io_out_valid(DFT2_bw32_24_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_25 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_25_clock),
    .reset(DFT2_bw32_25_reset),
    .io_in_en(DFT2_bw32_25_io_in_en),
    .io_in_valid(DFT2_bw32_25_io_in_valid),
    .io_in_0_Re(DFT2_bw32_25_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_25_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_25_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_25_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_25_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_25_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_25_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_25_io_out_1_Im),
    .io_out_valid(DFT2_bw32_25_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_26 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_26_clock),
    .reset(DFT2_bw32_26_reset),
    .io_in_en(DFT2_bw32_26_io_in_en),
    .io_in_valid(DFT2_bw32_26_io_in_valid),
    .io_in_0_Re(DFT2_bw32_26_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_26_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_26_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_26_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_26_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_26_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_26_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_26_io_out_1_Im),
    .io_out_valid(DFT2_bw32_26_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_27 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_27_clock),
    .reset(DFT2_bw32_27_reset),
    .io_in_en(DFT2_bw32_27_io_in_en),
    .io_in_valid(DFT2_bw32_27_io_in_valid),
    .io_in_0_Re(DFT2_bw32_27_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_27_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_27_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_27_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_27_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_27_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_27_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_27_io_out_1_Im),
    .io_out_valid(DFT2_bw32_27_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_28 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_28_clock),
    .reset(DFT2_bw32_28_reset),
    .io_in_en(DFT2_bw32_28_io_in_en),
    .io_in_valid(DFT2_bw32_28_io_in_valid),
    .io_in_0_Re(DFT2_bw32_28_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_28_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_28_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_28_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_28_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_28_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_28_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_28_io_out_1_Im),
    .io_out_valid(DFT2_bw32_28_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_29 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_29_clock),
    .reset(DFT2_bw32_29_reset),
    .io_in_en(DFT2_bw32_29_io_in_en),
    .io_in_valid(DFT2_bw32_29_io_in_valid),
    .io_in_0_Re(DFT2_bw32_29_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_29_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_29_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_29_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_29_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_29_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_29_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_29_io_out_1_Im),
    .io_out_valid(DFT2_bw32_29_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_30 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_30_clock),
    .reset(DFT2_bw32_30_reset),
    .io_in_en(DFT2_bw32_30_io_in_en),
    .io_in_valid(DFT2_bw32_30_io_in_valid),
    .io_in_0_Re(DFT2_bw32_30_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_30_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_30_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_30_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_30_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_30_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_30_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_30_io_out_1_Im),
    .io_out_valid(DFT2_bw32_30_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_31 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_31_clock),
    .reset(DFT2_bw32_31_reset),
    .io_in_en(DFT2_bw32_31_io_in_en),
    .io_in_valid(DFT2_bw32_31_io_in_valid),
    .io_in_0_Re(DFT2_bw32_31_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_31_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_31_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_31_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_31_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_31_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_31_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_31_io_out_1_Im),
    .io_out_valid(DFT2_bw32_31_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_32 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_32_clock),
    .reset(DFT2_bw32_32_reset),
    .io_in_en(DFT2_bw32_32_io_in_en),
    .io_in_valid(DFT2_bw32_32_io_in_valid),
    .io_in_0_Re(DFT2_bw32_32_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_32_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_32_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_32_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_32_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_32_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_32_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_32_io_out_1_Im),
    .io_out_valid(DFT2_bw32_32_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_33 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_33_clock),
    .reset(DFT2_bw32_33_reset),
    .io_in_en(DFT2_bw32_33_io_in_en),
    .io_in_valid(DFT2_bw32_33_io_in_valid),
    .io_in_0_Re(DFT2_bw32_33_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_33_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_33_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_33_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_33_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_33_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_33_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_33_io_out_1_Im),
    .io_out_valid(DFT2_bw32_33_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_34 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_34_clock),
    .reset(DFT2_bw32_34_reset),
    .io_in_en(DFT2_bw32_34_io_in_en),
    .io_in_valid(DFT2_bw32_34_io_in_valid),
    .io_in_0_Re(DFT2_bw32_34_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_34_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_34_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_34_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_34_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_34_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_34_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_34_io_out_1_Im),
    .io_out_valid(DFT2_bw32_34_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_35 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_35_clock),
    .reset(DFT2_bw32_35_reset),
    .io_in_en(DFT2_bw32_35_io_in_en),
    .io_in_valid(DFT2_bw32_35_io_in_valid),
    .io_in_0_Re(DFT2_bw32_35_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_35_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_35_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_35_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_35_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_35_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_35_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_35_io_out_1_Im),
    .io_out_valid(DFT2_bw32_35_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_36 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_36_clock),
    .reset(DFT2_bw32_36_reset),
    .io_in_en(DFT2_bw32_36_io_in_en),
    .io_in_valid(DFT2_bw32_36_io_in_valid),
    .io_in_0_Re(DFT2_bw32_36_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_36_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_36_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_36_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_36_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_36_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_36_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_36_io_out_1_Im),
    .io_out_valid(DFT2_bw32_36_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_37 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_37_clock),
    .reset(DFT2_bw32_37_reset),
    .io_in_en(DFT2_bw32_37_io_in_en),
    .io_in_valid(DFT2_bw32_37_io_in_valid),
    .io_in_0_Re(DFT2_bw32_37_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_37_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_37_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_37_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_37_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_37_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_37_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_37_io_out_1_Im),
    .io_out_valid(DFT2_bw32_37_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_38 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_38_clock),
    .reset(DFT2_bw32_38_reset),
    .io_in_en(DFT2_bw32_38_io_in_en),
    .io_in_valid(DFT2_bw32_38_io_in_valid),
    .io_in_0_Re(DFT2_bw32_38_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_38_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_38_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_38_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_38_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_38_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_38_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_38_io_out_1_Im),
    .io_out_valid(DFT2_bw32_38_io_out_valid)
  );
  DFT2_bw32 DFT2_bw32_39 ( // @[FFTSRDesigns.scala 79:70]
    .clock(DFT2_bw32_39_clock),
    .reset(DFT2_bw32_39_reset),
    .io_in_en(DFT2_bw32_39_io_in_en),
    .io_in_valid(DFT2_bw32_39_io_in_valid),
    .io_in_0_Re(DFT2_bw32_39_io_in_0_Re),
    .io_in_0_Im(DFT2_bw32_39_io_in_0_Im),
    .io_in_1_Re(DFT2_bw32_39_io_in_1_Re),
    .io_in_1_Im(DFT2_bw32_39_io_in_1_Im),
    .io_out_0_Re(DFT2_bw32_39_io_out_0_Re),
    .io_out_0_Im(DFT2_bw32_39_io_out_0_Im),
    .io_out_1_Re(DFT2_bw32_39_io_out_1_Re),
    .io_out_1_Im(DFT2_bw32_39_io_out_1_Im),
    .io_out_valid(DFT2_bw32_39_io_out_valid)
  );
  Permute_Streaming_N32_r2_w16_bitRtrue_bw64 Permute_Streaming_N32_r2_w16_bitRtrue_bw64 ( // @[FFTSRDesigns.scala 82:15]
    .clock(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_clock),
    .reset(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_reset),
    .io_in_en(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_en),
    .io_in_0(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_0),
    .io_in_1(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_1),
    .io_in_2(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_2),
    .io_in_3(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_3),
    .io_in_4(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_4),
    .io_in_5(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_5),
    .io_in_6(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_6),
    .io_in_7(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_7),
    .io_in_8(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_8),
    .io_in_9(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_9),
    .io_in_10(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_10),
    .io_in_11(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_11),
    .io_in_12(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_12),
    .io_in_13(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_13),
    .io_in_14(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_14),
    .io_in_15(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_15),
    .io_in_valid(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_valid),
    .io_out_0(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_0),
    .io_out_1(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_1),
    .io_out_2(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_2),
    .io_out_3(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_3),
    .io_out_4(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_4),
    .io_out_5(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_5),
    .io_out_6(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_6),
    .io_out_7(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_7),
    .io_out_8(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_8),
    .io_out_9(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_9),
    .io_out_10(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_10),
    .io_out_11(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_11),
    .io_out_12(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_12),
    .io_out_13(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_13),
    .io_out_14(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_14),
    .io_out_15(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_15),
    .io_out_valid(Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_valid)
  );
  Permute_Streaming_N32_r2_w16_bitRfalse_bw64 Permute_Streaming_N32_r2_w16_bitRfalse_bw64 ( // @[FFTSRDesigns.scala 84:15]
    .clock(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_clock),
    .reset(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_reset),
    .io_in_en(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_en),
    .io_in_0(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_0),
    .io_in_1(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_1),
    .io_in_2(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_2),
    .io_in_3(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_3),
    .io_in_4(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_4),
    .io_in_5(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_5),
    .io_in_6(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_6),
    .io_in_7(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_7),
    .io_in_8(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_8),
    .io_in_9(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_9),
    .io_in_10(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_10),
    .io_in_11(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_11),
    .io_in_12(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_12),
    .io_in_13(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_13),
    .io_in_14(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_14),
    .io_in_15(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_15),
    .io_in_valid(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_valid),
    .io_out_0(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_0),
    .io_out_1(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_1),
    .io_out_2(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_2),
    .io_out_3(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_3),
    .io_out_4(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_4),
    .io_out_5(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_5),
    .io_out_6(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_6),
    .io_out_7(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_7),
    .io_out_8(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_8),
    .io_out_9(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_9),
    .io_out_10(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_10),
    .io_out_11(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_11),
    .io_out_12(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_12),
    .io_out_13(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_13),
    .io_out_14(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_14),
    .io_out_15(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_15),
    .io_out_valid(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_valid)
  );
  Permute_Streaming_N32_r2_w16_bitRfalse_bw64 Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1 ( // @[FFTSRDesigns.scala 84:15]
    .clock(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_clock),
    .reset(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_reset),
    .io_in_en(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_en),
    .io_in_0(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_0),
    .io_in_1(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_1),
    .io_in_2(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_2),
    .io_in_3(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_3),
    .io_in_4(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_4),
    .io_in_5(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_5),
    .io_in_6(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_6),
    .io_in_7(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_7),
    .io_in_8(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_8),
    .io_in_9(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_9),
    .io_in_10(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_10),
    .io_in_11(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_11),
    .io_in_12(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_12),
    .io_in_13(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_13),
    .io_in_14(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_14),
    .io_in_15(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_15),
    .io_in_valid(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_valid),
    .io_out_0(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_0),
    .io_out_1(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_1),
    .io_out_2(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_2),
    .io_out_3(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_3),
    .io_out_4(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_4),
    .io_out_5(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_5),
    .io_out_6(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_6),
    .io_out_7(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_7),
    .io_out_8(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_8),
    .io_out_9(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_9),
    .io_out_10(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_10),
    .io_out_11(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_11),
    .io_out_12(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_12),
    .io_out_13(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_13),
    .io_out_14(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_14),
    .io_out_15(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_15),
    .io_out_valid(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_valid)
  );
  Permute_Streaming_N32_r2_w16_bitRfalse_bw64 Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2 ( // @[FFTSRDesigns.scala 84:15]
    .clock(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_clock),
    .reset(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_reset),
    .io_in_en(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_en),
    .io_in_0(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_0),
    .io_in_1(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_1),
    .io_in_2(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_2),
    .io_in_3(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_3),
    .io_in_4(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_4),
    .io_in_5(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_5),
    .io_in_6(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_6),
    .io_in_7(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_7),
    .io_in_8(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_8),
    .io_in_9(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_9),
    .io_in_10(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_10),
    .io_in_11(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_11),
    .io_in_12(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_12),
    .io_in_13(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_13),
    .io_in_14(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_14),
    .io_in_15(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_15),
    .io_in_valid(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_valid),
    .io_out_0(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_0),
    .io_out_1(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_1),
    .io_out_2(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_2),
    .io_out_3(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_3),
    .io_out_4(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_4),
    .io_out_5(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_5),
    .io_out_6(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_6),
    .io_out_7(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_7),
    .io_out_8(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_8),
    .io_out_9(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_9),
    .io_out_10(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_10),
    .io_out_11(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_11),
    .io_out_12(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_12),
    .io_out_13(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_13),
    .io_out_14(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_14),
    .io_out_15(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_15),
    .io_out_valid(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_valid)
  );
  Permute_Streaming_N32_r2_w16_bitRfalse_bw64 Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3 ( // @[FFTSRDesigns.scala 84:15]
    .clock(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_clock),
    .reset(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_reset),
    .io_in_en(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_en),
    .io_in_0(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_0),
    .io_in_1(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_1),
    .io_in_2(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_2),
    .io_in_3(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_3),
    .io_in_4(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_4),
    .io_in_5(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_5),
    .io_in_6(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_6),
    .io_in_7(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_7),
    .io_in_8(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_8),
    .io_in_9(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_9),
    .io_in_10(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_10),
    .io_in_11(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_11),
    .io_in_12(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_12),
    .io_in_13(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_13),
    .io_in_14(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_14),
    .io_in_15(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_15),
    .io_in_valid(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_valid),
    .io_out_0(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_0),
    .io_out_1(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_1),
    .io_out_2(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_2),
    .io_out_3(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_3),
    .io_out_4(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_4),
    .io_out_5(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_5),
    .io_out_6(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_6),
    .io_out_7(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_7),
    .io_out_8(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_8),
    .io_out_9(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_9),
    .io_out_10(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_10),
    .io_out_11(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_11),
    .io_out_12(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_12),
    .io_out_13(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_13),
    .io_out_14(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_14),
    .io_out_15(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_15),
    .io_out_valid(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_valid)
  );
  Permute_Streaming_N32_r2_w16_bitRfalse_bw64 Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4 ( // @[FFTSRDesigns.scala 84:15]
    .clock(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_clock),
    .reset(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_reset),
    .io_in_en(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_en),
    .io_in_0(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_0),
    .io_in_1(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_1),
    .io_in_2(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_2),
    .io_in_3(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_3),
    .io_in_4(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_4),
    .io_in_5(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_5),
    .io_in_6(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_6),
    .io_in_7(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_7),
    .io_in_8(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_8),
    .io_in_9(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_9),
    .io_in_10(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_10),
    .io_in_11(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_11),
    .io_in_12(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_12),
    .io_in_13(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_13),
    .io_in_14(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_14),
    .io_in_15(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_15),
    .io_in_valid(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_valid),
    .io_out_0(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_0),
    .io_out_1(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_1),
    .io_out_2(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_2),
    .io_out_3(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_3),
    .io_out_4(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_4),
    .io_out_5(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_5),
    .io_out_6(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_6),
    .io_out_7(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_7),
    .io_out_8(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_8),
    .io_out_9(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_9),
    .io_out_10(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_10),
    .io_out_11(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_11),
    .io_out_12(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_12),
    .io_out_13(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_13),
    .io_out_14(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_14),
    .io_out_15(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_15),
    .io_out_valid(Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_valid)
  );
  TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32 TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32 ( // @[FFTSRDesigns.scala 86:68]
    .clock(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_clock),
    .reset(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_reset),
    .io_in_inv(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_inv),
    .io_in_en(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_en),
    .io_in_0_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_0_Re),
    .io_in_0_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_0_Im),
    .io_in_1_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_1_Re),
    .io_in_1_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_1_Im),
    .io_in_2_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_2_Re),
    .io_in_2_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_2_Im),
    .io_in_3_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_3_Re),
    .io_in_3_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_3_Im),
    .io_in_4_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_4_Re),
    .io_in_4_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_4_Im),
    .io_in_5_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_5_Re),
    .io_in_5_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_5_Im),
    .io_in_6_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_6_Re),
    .io_in_6_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_6_Im),
    .io_in_7_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_7_Re),
    .io_in_7_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_7_Im),
    .io_in_8_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_8_Re),
    .io_in_8_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_8_Im),
    .io_in_9_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_9_Re),
    .io_in_9_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_9_Im),
    .io_in_10_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_10_Re),
    .io_in_10_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_10_Im),
    .io_in_11_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_11_Re),
    .io_in_11_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_11_Im),
    .io_in_12_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_12_Re),
    .io_in_12_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_12_Im),
    .io_in_13_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_13_Re),
    .io_in_13_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_13_Im),
    .io_in_14_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_14_Re),
    .io_in_14_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_14_Im),
    .io_in_15_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_15_Re),
    .io_in_15_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_15_Im),
    .io_in_valid(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_valid),
    .io_out_valid(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_valid),
    .io_out_0_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_0_Re),
    .io_out_0_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_0_Im),
    .io_out_1_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_1_Re),
    .io_out_1_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_1_Im),
    .io_out_2_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_2_Re),
    .io_out_2_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_2_Im),
    .io_out_3_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_3_Re),
    .io_out_3_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_3_Im),
    .io_out_4_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_4_Re),
    .io_out_4_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_4_Im),
    .io_out_5_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_5_Re),
    .io_out_5_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_5_Im),
    .io_out_6_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_6_Re),
    .io_out_6_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_6_Im),
    .io_out_7_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_7_Re),
    .io_out_7_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_7_Im),
    .io_out_8_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_8_Re),
    .io_out_8_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_8_Im),
    .io_out_9_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_9_Re),
    .io_out_9_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_9_Im),
    .io_out_10_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_10_Re),
    .io_out_10_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_10_Im),
    .io_out_11_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_11_Re),
    .io_out_11_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_11_Im),
    .io_out_12_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_12_Re),
    .io_out_12_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_12_Im),
    .io_out_13_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_13_Re),
    .io_out_13_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_13_Im),
    .io_out_14_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_14_Re),
    .io_out_14_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_14_Im),
    .io_out_15_Re(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_15_Re),
    .io_out_15_Im(TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_15_Im)
  );
  TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32 TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32 ( // @[FFTSRDesigns.scala 86:68]
    .clock(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_clock),
    .reset(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_reset),
    .io_in_inv(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_inv),
    .io_in_en(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_en),
    .io_in_0_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_0_Re),
    .io_in_0_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_0_Im),
    .io_in_1_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_1_Re),
    .io_in_1_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_1_Im),
    .io_in_2_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_2_Re),
    .io_in_2_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_2_Im),
    .io_in_3_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_3_Re),
    .io_in_3_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_3_Im),
    .io_in_4_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_4_Re),
    .io_in_4_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_4_Im),
    .io_in_5_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_5_Re),
    .io_in_5_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_5_Im),
    .io_in_6_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_6_Re),
    .io_in_6_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_6_Im),
    .io_in_7_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_7_Re),
    .io_in_7_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_7_Im),
    .io_in_8_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_8_Re),
    .io_in_8_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_8_Im),
    .io_in_9_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_9_Re),
    .io_in_9_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_9_Im),
    .io_in_10_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_10_Re),
    .io_in_10_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_10_Im),
    .io_in_11_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_11_Re),
    .io_in_11_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_11_Im),
    .io_in_12_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_12_Re),
    .io_in_12_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_12_Im),
    .io_in_13_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_13_Re),
    .io_in_13_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_13_Im),
    .io_in_14_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_14_Re),
    .io_in_14_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_14_Im),
    .io_in_15_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_15_Re),
    .io_in_15_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_15_Im),
    .io_in_valid(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_valid),
    .io_out_valid(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_valid),
    .io_out_0_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_0_Re),
    .io_out_0_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_0_Im),
    .io_out_1_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_1_Re),
    .io_out_1_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_1_Im),
    .io_out_2_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_2_Re),
    .io_out_2_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_2_Im),
    .io_out_3_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_3_Re),
    .io_out_3_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_3_Im),
    .io_out_4_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_4_Re),
    .io_out_4_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_4_Im),
    .io_out_5_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_5_Re),
    .io_out_5_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_5_Im),
    .io_out_6_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_6_Re),
    .io_out_6_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_6_Im),
    .io_out_7_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_7_Re),
    .io_out_7_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_7_Im),
    .io_out_8_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_8_Re),
    .io_out_8_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_8_Im),
    .io_out_9_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_9_Re),
    .io_out_9_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_9_Im),
    .io_out_10_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_10_Re),
    .io_out_10_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_10_Im),
    .io_out_11_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_11_Re),
    .io_out_11_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_11_Im),
    .io_out_12_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_12_Re),
    .io_out_12_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_12_Im),
    .io_out_13_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_13_Re),
    .io_out_13_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_13_Im),
    .io_out_14_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_14_Re),
    .io_out_14_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_14_Im),
    .io_out_15_Re(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_15_Re),
    .io_out_15_Im(TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_15_Im)
  );
  TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32 TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32 ( // @[FFTSRDesigns.scala 86:68]
    .clock(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_clock),
    .reset(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_reset),
    .io_in_inv(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_inv),
    .io_in_en(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_en),
    .io_in_0_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_0_Re),
    .io_in_0_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_0_Im),
    .io_in_1_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_1_Re),
    .io_in_1_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_1_Im),
    .io_in_2_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_2_Re),
    .io_in_2_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_2_Im),
    .io_in_3_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_3_Re),
    .io_in_3_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_3_Im),
    .io_in_4_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_4_Re),
    .io_in_4_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_4_Im),
    .io_in_5_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_5_Re),
    .io_in_5_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_5_Im),
    .io_in_6_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_6_Re),
    .io_in_6_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_6_Im),
    .io_in_7_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_7_Re),
    .io_in_7_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_7_Im),
    .io_in_8_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_8_Re),
    .io_in_8_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_8_Im),
    .io_in_9_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_9_Re),
    .io_in_9_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_9_Im),
    .io_in_10_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_10_Re),
    .io_in_10_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_10_Im),
    .io_in_11_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_11_Re),
    .io_in_11_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_11_Im),
    .io_in_12_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_12_Re),
    .io_in_12_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_12_Im),
    .io_in_13_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_13_Re),
    .io_in_13_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_13_Im),
    .io_in_14_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_14_Re),
    .io_in_14_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_14_Im),
    .io_in_15_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_15_Re),
    .io_in_15_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_15_Im),
    .io_in_valid(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_valid),
    .io_out_valid(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_valid),
    .io_out_0_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_0_Re),
    .io_out_0_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_0_Im),
    .io_out_1_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_1_Re),
    .io_out_1_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_1_Im),
    .io_out_2_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_2_Re),
    .io_out_2_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_2_Im),
    .io_out_3_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_3_Re),
    .io_out_3_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_3_Im),
    .io_out_4_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_4_Re),
    .io_out_4_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_4_Im),
    .io_out_5_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_5_Re),
    .io_out_5_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_5_Im),
    .io_out_6_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_6_Re),
    .io_out_6_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_6_Im),
    .io_out_7_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_7_Re),
    .io_out_7_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_7_Im),
    .io_out_8_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_8_Re),
    .io_out_8_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_8_Im),
    .io_out_9_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_9_Re),
    .io_out_9_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_9_Im),
    .io_out_10_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_10_Re),
    .io_out_10_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_10_Im),
    .io_out_11_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_11_Re),
    .io_out_11_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_11_Im),
    .io_out_12_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_12_Re),
    .io_out_12_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_12_Im),
    .io_out_13_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_13_Re),
    .io_out_13_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_13_Im),
    .io_out_14_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_14_Re),
    .io_out_14_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_14_Im),
    .io_out_15_Re(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_15_Re),
    .io_out_15_Im(TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_15_Im)
  );
  TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32 TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32 ( // @[FFTSRDesigns.scala 86:68]
    .clock(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_clock),
    .reset(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_reset),
    .io_in_inv(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_inv),
    .io_in_en(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_en),
    .io_in_0_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_0_Re),
    .io_in_0_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_0_Im),
    .io_in_1_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_1_Re),
    .io_in_1_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_1_Im),
    .io_in_2_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_2_Re),
    .io_in_2_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_2_Im),
    .io_in_3_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_3_Re),
    .io_in_3_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_3_Im),
    .io_in_4_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_4_Re),
    .io_in_4_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_4_Im),
    .io_in_5_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_5_Re),
    .io_in_5_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_5_Im),
    .io_in_6_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_6_Re),
    .io_in_6_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_6_Im),
    .io_in_7_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_7_Re),
    .io_in_7_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_7_Im),
    .io_in_8_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_8_Re),
    .io_in_8_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_8_Im),
    .io_in_9_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_9_Re),
    .io_in_9_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_9_Im),
    .io_in_10_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_10_Re),
    .io_in_10_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_10_Im),
    .io_in_11_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_11_Re),
    .io_in_11_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_11_Im),
    .io_in_12_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_12_Re),
    .io_in_12_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_12_Im),
    .io_in_13_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_13_Re),
    .io_in_13_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_13_Im),
    .io_in_14_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_14_Re),
    .io_in_14_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_14_Im),
    .io_in_15_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_15_Re),
    .io_in_15_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_15_Im),
    .io_in_valid(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_valid),
    .io_out_valid(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_valid),
    .io_out_0_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_0_Re),
    .io_out_0_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_0_Im),
    .io_out_1_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_1_Re),
    .io_out_1_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_1_Im),
    .io_out_2_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_2_Re),
    .io_out_2_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_2_Im),
    .io_out_3_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_3_Re),
    .io_out_3_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_3_Im),
    .io_out_4_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_4_Re),
    .io_out_4_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_4_Im),
    .io_out_5_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_5_Re),
    .io_out_5_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_5_Im),
    .io_out_6_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_6_Re),
    .io_out_6_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_6_Im),
    .io_out_7_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_7_Re),
    .io_out_7_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_7_Im),
    .io_out_8_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_8_Re),
    .io_out_8_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_8_Im),
    .io_out_9_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_9_Re),
    .io_out_9_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_9_Im),
    .io_out_10_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_10_Re),
    .io_out_10_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_10_Im),
    .io_out_11_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_11_Re),
    .io_out_11_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_11_Im),
    .io_out_12_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_12_Re),
    .io_out_12_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_12_Im),
    .io_out_13_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_13_Re),
    .io_out_13_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_13_Im),
    .io_out_14_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_14_Re),
    .io_out_14_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_14_Im),
    .io_out_15_Re(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_15_Re),
    .io_out_15_Im(TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_15_Im)
  );
  assign io_out_valid = Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_out_valid; // @[FFTSRDesigns.scala 88:18]
  assign io_out_0_Re = _WIRE_1[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_0_Im = _WIRE_1[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_1_Re = _WIRE_3[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_1_Im = _WIRE_3[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_2_Re = _WIRE_5[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_2_Im = _WIRE_5[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_3_Re = _WIRE_7[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_3_Im = _WIRE_7[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_4_Re = _WIRE_9[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_4_Im = _WIRE_9[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_5_Re = _WIRE_11[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_5_Im = _WIRE_11[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_6_Re = _WIRE_13[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_6_Im = _WIRE_13[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_7_Re = _WIRE_15[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_7_Im = _WIRE_15[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_8_Re = _WIRE_17[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_8_Im = _WIRE_17[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_9_Re = _WIRE_19[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_9_Im = _WIRE_19[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_10_Re = _WIRE_21[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_10_Im = _WIRE_21[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_11_Re = _WIRE_23[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_11_Im = _WIRE_23[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_12_Re = _WIRE_25[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_12_Im = _WIRE_25[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_13_Re = _WIRE_27[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_13_Im = _WIRE_27[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_14_Re = _WIRE_29[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_14_Im = _WIRE_29[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_15_Re = _WIRE_31[63:32]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_15_Im = _WIRE_31[31:0]; // @[FFTSRDesigns.scala 89:72]
  assign io_out_ready = io_in_ready; // @[FFTSRDesigns.scala 87:18]
  assign DFT2_bw32_clock = clock;
  assign DFT2_bw32_reset = reset;
  assign DFT2_bw32_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_io_in_valid = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_valid; // @[FFTSRDesigns.scala 108:38]
  assign DFT2_bw32_io_in_0_Re = _WIRE_44[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_io_in_0_Im = _WIRE_44[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_io_in_1_Re = _WIRE_46[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_io_in_1_Im = _WIRE_46[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_1_clock = clock;
  assign DFT2_bw32_1_reset = reset;
  assign DFT2_bw32_1_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_1_io_in_valid = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_valid; // @[FFTSRDesigns.scala 108:38]
  assign DFT2_bw32_1_io_in_0_Re = _WIRE_49[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_1_io_in_0_Im = _WIRE_49[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_1_io_in_1_Re = _WIRE_51[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_1_io_in_1_Im = _WIRE_51[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_2_clock = clock;
  assign DFT2_bw32_2_reset = reset;
  assign DFT2_bw32_2_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_2_io_in_valid = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_valid; // @[FFTSRDesigns.scala 108:38]
  assign DFT2_bw32_2_io_in_0_Re = _WIRE_54[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_2_io_in_0_Im = _WIRE_54[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_2_io_in_1_Re = _WIRE_56[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_2_io_in_1_Im = _WIRE_56[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_3_clock = clock;
  assign DFT2_bw32_3_reset = reset;
  assign DFT2_bw32_3_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_3_io_in_valid = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_valid; // @[FFTSRDesigns.scala 108:38]
  assign DFT2_bw32_3_io_in_0_Re = _WIRE_59[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_3_io_in_0_Im = _WIRE_59[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_3_io_in_1_Re = _WIRE_61[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_3_io_in_1_Im = _WIRE_61[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_4_clock = clock;
  assign DFT2_bw32_4_reset = reset;
  assign DFT2_bw32_4_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_4_io_in_valid = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_valid; // @[FFTSRDesigns.scala 108:38]
  assign DFT2_bw32_4_io_in_0_Re = _WIRE_64[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_4_io_in_0_Im = _WIRE_64[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_4_io_in_1_Re = _WIRE_66[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_4_io_in_1_Im = _WIRE_66[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_5_clock = clock;
  assign DFT2_bw32_5_reset = reset;
  assign DFT2_bw32_5_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_5_io_in_valid = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_valid; // @[FFTSRDesigns.scala 108:38]
  assign DFT2_bw32_5_io_in_0_Re = _WIRE_69[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_5_io_in_0_Im = _WIRE_69[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_5_io_in_1_Re = _WIRE_71[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_5_io_in_1_Im = _WIRE_71[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_6_clock = clock;
  assign DFT2_bw32_6_reset = reset;
  assign DFT2_bw32_6_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_6_io_in_valid = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_valid; // @[FFTSRDesigns.scala 108:38]
  assign DFT2_bw32_6_io_in_0_Re = _WIRE_74[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_6_io_in_0_Im = _WIRE_74[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_6_io_in_1_Re = _WIRE_76[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_6_io_in_1_Im = _WIRE_76[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_7_clock = clock;
  assign DFT2_bw32_7_reset = reset;
  assign DFT2_bw32_7_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_7_io_in_valid = Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_out_valid; // @[FFTSRDesigns.scala 108:38]
  assign DFT2_bw32_7_io_in_0_Re = _WIRE_79[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_7_io_in_0_Im = _WIRE_79[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_7_io_in_1_Re = _WIRE_81[63:32]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_7_io_in_1_Im = _WIRE_81[31:0]; // @[FFTSRDesigns.scala 109:96]
  assign DFT2_bw32_8_clock = clock;
  assign DFT2_bw32_8_reset = reset;
  assign DFT2_bw32_8_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_8_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_8_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_0_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_8_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_0_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_8_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_1_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_8_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_1_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_9_clock = clock;
  assign DFT2_bw32_9_reset = reset;
  assign DFT2_bw32_9_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_9_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_9_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_2_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_9_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_2_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_9_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_3_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_9_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_3_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_10_clock = clock;
  assign DFT2_bw32_10_reset = reset;
  assign DFT2_bw32_10_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_10_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_10_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_4_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_10_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_4_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_10_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_5_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_10_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_5_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_11_clock = clock;
  assign DFT2_bw32_11_reset = reset;
  assign DFT2_bw32_11_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_11_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_11_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_6_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_11_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_6_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_11_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_7_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_11_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_7_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_12_clock = clock;
  assign DFT2_bw32_12_reset = reset;
  assign DFT2_bw32_12_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_12_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_12_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_8_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_12_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_8_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_12_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_9_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_12_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_9_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_13_clock = clock;
  assign DFT2_bw32_13_reset = reset;
  assign DFT2_bw32_13_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_13_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_13_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_10_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_13_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_10_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_13_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_11_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_13_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_11_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_14_clock = clock;
  assign DFT2_bw32_14_reset = reset;
  assign DFT2_bw32_14_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_14_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_14_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_12_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_14_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_12_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_14_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_13_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_14_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_13_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_15_clock = clock;
  assign DFT2_bw32_15_reset = reset;
  assign DFT2_bw32_15_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_15_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_15_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_14_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_15_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_14_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_15_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_15_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_15_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_out_15_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_16_clock = clock;
  assign DFT2_bw32_16_reset = reset;
  assign DFT2_bw32_16_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_16_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_16_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_0_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_16_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_0_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_16_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_1_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_16_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_1_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_17_clock = clock;
  assign DFT2_bw32_17_reset = reset;
  assign DFT2_bw32_17_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_17_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_17_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_2_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_17_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_2_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_17_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_3_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_17_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_3_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_18_clock = clock;
  assign DFT2_bw32_18_reset = reset;
  assign DFT2_bw32_18_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_18_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_18_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_4_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_18_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_4_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_18_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_5_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_18_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_5_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_19_clock = clock;
  assign DFT2_bw32_19_reset = reset;
  assign DFT2_bw32_19_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_19_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_19_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_6_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_19_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_6_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_19_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_7_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_19_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_7_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_20_clock = clock;
  assign DFT2_bw32_20_reset = reset;
  assign DFT2_bw32_20_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_20_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_20_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_8_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_20_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_8_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_20_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_9_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_20_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_9_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_21_clock = clock;
  assign DFT2_bw32_21_reset = reset;
  assign DFT2_bw32_21_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_21_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_21_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_10_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_21_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_10_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_21_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_11_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_21_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_11_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_22_clock = clock;
  assign DFT2_bw32_22_reset = reset;
  assign DFT2_bw32_22_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_22_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_22_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_12_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_22_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_12_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_22_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_13_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_22_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_13_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_23_clock = clock;
  assign DFT2_bw32_23_reset = reset;
  assign DFT2_bw32_23_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_23_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_23_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_14_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_23_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_14_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_23_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_15_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_23_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_out_15_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_24_clock = clock;
  assign DFT2_bw32_24_reset = reset;
  assign DFT2_bw32_24_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_24_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_24_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_0_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_24_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_0_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_24_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_1_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_24_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_1_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_25_clock = clock;
  assign DFT2_bw32_25_reset = reset;
  assign DFT2_bw32_25_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_25_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_25_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_2_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_25_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_2_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_25_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_3_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_25_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_3_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_26_clock = clock;
  assign DFT2_bw32_26_reset = reset;
  assign DFT2_bw32_26_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_26_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_26_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_4_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_26_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_4_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_26_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_5_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_26_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_5_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_27_clock = clock;
  assign DFT2_bw32_27_reset = reset;
  assign DFT2_bw32_27_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_27_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_27_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_6_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_27_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_6_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_27_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_7_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_27_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_7_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_28_clock = clock;
  assign DFT2_bw32_28_reset = reset;
  assign DFT2_bw32_28_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_28_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_28_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_8_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_28_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_8_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_28_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_9_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_28_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_9_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_29_clock = clock;
  assign DFT2_bw32_29_reset = reset;
  assign DFT2_bw32_29_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_29_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_29_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_10_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_29_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_10_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_29_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_11_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_29_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_11_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_30_clock = clock;
  assign DFT2_bw32_30_reset = reset;
  assign DFT2_bw32_30_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_30_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_30_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_12_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_30_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_12_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_30_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_13_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_30_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_13_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_31_clock = clock;
  assign DFT2_bw32_31_reset = reset;
  assign DFT2_bw32_31_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_31_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_31_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_14_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_31_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_14_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_31_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_15_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_31_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_out_15_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_32_clock = clock;
  assign DFT2_bw32_32_reset = reset;
  assign DFT2_bw32_32_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_32_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_32_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_0_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_32_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_0_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_32_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_1_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_32_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_1_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_33_clock = clock;
  assign DFT2_bw32_33_reset = reset;
  assign DFT2_bw32_33_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_33_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_33_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_2_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_33_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_2_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_33_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_3_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_33_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_3_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_34_clock = clock;
  assign DFT2_bw32_34_reset = reset;
  assign DFT2_bw32_34_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_34_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_34_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_4_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_34_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_4_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_34_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_5_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_34_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_5_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_35_clock = clock;
  assign DFT2_bw32_35_reset = reset;
  assign DFT2_bw32_35_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_35_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_35_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_6_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_35_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_6_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_35_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_7_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_35_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_7_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_36_clock = clock;
  assign DFT2_bw32_36_reset = reset;
  assign DFT2_bw32_36_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_36_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_36_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_8_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_36_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_8_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_36_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_9_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_36_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_9_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_37_clock = clock;
  assign DFT2_bw32_37_reset = reset;
  assign DFT2_bw32_37_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_37_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_37_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_10_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_37_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_10_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_37_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_11_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_37_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_11_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_38_clock = clock;
  assign DFT2_bw32_38_reset = reset;
  assign DFT2_bw32_38_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_38_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_38_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_12_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_38_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_12_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_38_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_13_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_38_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_13_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_39_clock = clock;
  assign DFT2_bw32_39_reset = reset;
  assign DFT2_bw32_39_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 91:43]
  assign DFT2_bw32_39_io_in_valid = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_valid; // @[FFTSRDesigns.scala 111:38]
  assign DFT2_bw32_39_io_in_0_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_14_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_39_io_in_0_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_14_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_39_io_in_1_Re = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_15_Re; // @[FFTSRDesigns.scala 112:{42,42}]
  assign DFT2_bw32_39_io_in_1_Im = TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_out_15_Im; // @[FFTSRDesigns.scala 112:{42,42}]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_clock = clock;
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_reset = reset;
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 90:34]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_0 = {io_in_0_Re,io_in_0_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_1 = {io_in_1_Re,io_in_1_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_2 = {io_in_2_Re,io_in_2_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_3 = {io_in_3_Re,io_in_3_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_4 = {io_in_4_Re,io_in_4_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_5 = {io_in_5_Re,io_in_5_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_6 = {io_in_6_Re,io_in_6_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_7 = {io_in_7_Re,io_in_7_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_8 = {io_in_8_Re,io_in_8_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_9 = {io_in_9_Re,io_in_9_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_10 = {io_in_10_Re,io_in_10_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_11 = {io_in_11_Re,io_in_11_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_12 = {io_in_12_Re,io_in_12_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_13 = {io_in_13_Re,io_in_13_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_14 = {io_in_14_Re,io_in_14_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_15 = {io_in_15_Re,io_in_15_Im}; // @[FFTSRDesigns.scala 93:47]
  assign Permute_Streaming_N32_r2_w16_bitRtrue_bw64_io_in_valid = io_in_valid; // @[FFTSRDesigns.scala 94:30]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_clock = clock;
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_reset = reset;
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 90:34]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_0 = {DFT2_bw32_io_out_0_Re,DFT2_bw32_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_1 = {DFT2_bw32_io_out_1_Re,DFT2_bw32_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_2 = {DFT2_bw32_1_io_out_0_Re,DFT2_bw32_1_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_3 = {DFT2_bw32_1_io_out_1_Re,DFT2_bw32_1_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_4 = {DFT2_bw32_2_io_out_0_Re,DFT2_bw32_2_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_5 = {DFT2_bw32_2_io_out_1_Re,DFT2_bw32_2_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_6 = {DFT2_bw32_3_io_out_0_Re,DFT2_bw32_3_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_7 = {DFT2_bw32_3_io_out_1_Re,DFT2_bw32_3_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_8 = {DFT2_bw32_4_io_out_0_Re,DFT2_bw32_4_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_9 = {DFT2_bw32_4_io_out_1_Re,DFT2_bw32_4_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_10 = {DFT2_bw32_5_io_out_0_Re,DFT2_bw32_5_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_11 = {DFT2_bw32_5_io_out_1_Re,DFT2_bw32_5_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_12 = {DFT2_bw32_6_io_out_0_Re,DFT2_bw32_6_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_13 = {DFT2_bw32_6_io_out_1_Re,DFT2_bw32_6_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_14 = {DFT2_bw32_7_io_out_0_Re,DFT2_bw32_7_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_15 = {DFT2_bw32_7_io_out_1_Re,DFT2_bw32_7_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_in_valid = DFT2_bw32_io_out_valid; // @[FFTSRDesigns.scala 96:34]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_clock = clock;
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_reset = reset;
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 90:34]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_0 = {DFT2_bw32_8_io_out_0_Re,DFT2_bw32_8_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_1 = {DFT2_bw32_8_io_out_1_Re,DFT2_bw32_8_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_2 = {DFT2_bw32_9_io_out_0_Re,DFT2_bw32_9_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_3 = {DFT2_bw32_9_io_out_1_Re,DFT2_bw32_9_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_4 = {DFT2_bw32_10_io_out_0_Re,DFT2_bw32_10_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_5 = {DFT2_bw32_10_io_out_1_Re,DFT2_bw32_10_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_6 = {DFT2_bw32_11_io_out_0_Re,DFT2_bw32_11_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_7 = {DFT2_bw32_11_io_out_1_Re,DFT2_bw32_11_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_8 = {DFT2_bw32_12_io_out_0_Re,DFT2_bw32_12_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_9 = {DFT2_bw32_12_io_out_1_Re,DFT2_bw32_12_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_10 = {DFT2_bw32_13_io_out_0_Re,DFT2_bw32_13_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_11 = {DFT2_bw32_13_io_out_1_Re,DFT2_bw32_13_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_12 = {DFT2_bw32_14_io_out_0_Re,DFT2_bw32_14_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_13 = {DFT2_bw32_14_io_out_1_Re,DFT2_bw32_14_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_14 = {DFT2_bw32_15_io_out_0_Re,DFT2_bw32_15_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_15 = {DFT2_bw32_15_io_out_1_Re,DFT2_bw32_15_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_in_valid = DFT2_bw32_8_io_out_valid; // @[FFTSRDesigns.scala 96:34]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_clock = clock;
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_reset = reset;
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 90:34]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_0 = {DFT2_bw32_16_io_out_0_Re,DFT2_bw32_16_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_1 = {DFT2_bw32_16_io_out_1_Re,DFT2_bw32_16_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_2 = {DFT2_bw32_17_io_out_0_Re,DFT2_bw32_17_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_3 = {DFT2_bw32_17_io_out_1_Re,DFT2_bw32_17_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_4 = {DFT2_bw32_18_io_out_0_Re,DFT2_bw32_18_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_5 = {DFT2_bw32_18_io_out_1_Re,DFT2_bw32_18_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_6 = {DFT2_bw32_19_io_out_0_Re,DFT2_bw32_19_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_7 = {DFT2_bw32_19_io_out_1_Re,DFT2_bw32_19_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_8 = {DFT2_bw32_20_io_out_0_Re,DFT2_bw32_20_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_9 = {DFT2_bw32_20_io_out_1_Re,DFT2_bw32_20_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_10 = {DFT2_bw32_21_io_out_0_Re,DFT2_bw32_21_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_11 = {DFT2_bw32_21_io_out_1_Re,DFT2_bw32_21_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_12 = {DFT2_bw32_22_io_out_0_Re,DFT2_bw32_22_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_13 = {DFT2_bw32_22_io_out_1_Re,DFT2_bw32_22_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_14 = {DFT2_bw32_23_io_out_0_Re,DFT2_bw32_23_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_15 = {DFT2_bw32_23_io_out_1_Re,DFT2_bw32_23_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_in_valid = DFT2_bw32_16_io_out_valid; // @[FFTSRDesigns.scala 96:34]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_clock = clock;
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_reset = reset;
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 90:34]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_0 = {DFT2_bw32_24_io_out_0_Re,DFT2_bw32_24_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_1 = {DFT2_bw32_24_io_out_1_Re,DFT2_bw32_24_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_2 = {DFT2_bw32_25_io_out_0_Re,DFT2_bw32_25_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_3 = {DFT2_bw32_25_io_out_1_Re,DFT2_bw32_25_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_4 = {DFT2_bw32_26_io_out_0_Re,DFT2_bw32_26_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_5 = {DFT2_bw32_26_io_out_1_Re,DFT2_bw32_26_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_6 = {DFT2_bw32_27_io_out_0_Re,DFT2_bw32_27_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_7 = {DFT2_bw32_27_io_out_1_Re,DFT2_bw32_27_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_8 = {DFT2_bw32_28_io_out_0_Re,DFT2_bw32_28_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_9 = {DFT2_bw32_28_io_out_1_Re,DFT2_bw32_28_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_10 = {DFT2_bw32_29_io_out_0_Re,DFT2_bw32_29_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_11 = {DFT2_bw32_29_io_out_1_Re,DFT2_bw32_29_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_12 = {DFT2_bw32_30_io_out_0_Re,DFT2_bw32_30_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_13 = {DFT2_bw32_30_io_out_1_Re,DFT2_bw32_30_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_14 = {DFT2_bw32_31_io_out_0_Re,DFT2_bw32_31_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_15 = {DFT2_bw32_31_io_out_1_Re,DFT2_bw32_31_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_in_valid = DFT2_bw32_24_io_out_valid; // @[FFTSRDesigns.scala 96:34]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_clock = clock;
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_reset = reset;
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 90:34]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_0 = {DFT2_bw32_32_io_out_0_Re,DFT2_bw32_32_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_1 = {DFT2_bw32_32_io_out_1_Re,DFT2_bw32_32_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_2 = {DFT2_bw32_33_io_out_0_Re,DFT2_bw32_33_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_3 = {DFT2_bw32_33_io_out_1_Re,DFT2_bw32_33_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_4 = {DFT2_bw32_34_io_out_0_Re,DFT2_bw32_34_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_5 = {DFT2_bw32_34_io_out_1_Re,DFT2_bw32_34_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_6 = {DFT2_bw32_35_io_out_0_Re,DFT2_bw32_35_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_7 = {DFT2_bw32_35_io_out_1_Re,DFT2_bw32_35_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_8 = {DFT2_bw32_36_io_out_0_Re,DFT2_bw32_36_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_9 = {DFT2_bw32_36_io_out_1_Re,DFT2_bw32_36_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_10 = {DFT2_bw32_37_io_out_0_Re,DFT2_bw32_37_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_11 = {DFT2_bw32_37_io_out_1_Re,DFT2_bw32_37_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_12 = {DFT2_bw32_38_io_out_0_Re,DFT2_bw32_38_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_13 = {DFT2_bw32_38_io_out_1_Re,DFT2_bw32_38_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_14 = {DFT2_bw32_39_io_out_0_Re,DFT2_bw32_39_io_out_0_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_15 = {DFT2_bw32_39_io_out_1_Re,DFT2_bw32_39_io_out_1_Im}; // @[FFTSRDesigns.scala 98:45]
  assign Permute_Streaming_N32_r2_w16_bitRfalse_bw64_4_io_in_valid = DFT2_bw32_32_io_out_valid; // @[FFTSRDesigns.scala 96:34]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_clock = clock;
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_reset = reset;
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_inv = io_in_inv; // @[FFTSRDesigns.scala 101:34]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 92:34]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_0_Re = _WIRE_93[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_0_Im = _WIRE_93[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_1_Re = _WIRE_95[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_1_Im = _WIRE_95[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_2_Re = _WIRE_97[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_2_Im = _WIRE_97[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_3_Re = _WIRE_99[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_3_Im = _WIRE_99[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_4_Re = _WIRE_101[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_4_Im = _WIRE_101[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_5_Re = _WIRE_103[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_5_Im = _WIRE_103[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_6_Re = _WIRE_105[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_6_Im = _WIRE_105[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_7_Re = _WIRE_107[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_7_Im = _WIRE_107[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_8_Re = _WIRE_109[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_8_Im = _WIRE_109[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_9_Re = _WIRE_111[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_9_Im = _WIRE_111[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_10_Re = _WIRE_113[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_10_Im = _WIRE_113[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_11_Re = _WIRE_115[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_11_Im = _WIRE_115[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_12_Re = _WIRE_117[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_12_Im = _WIRE_117[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_13_Re = _WIRE_119[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_13_Im = _WIRE_119[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_14_Re = _WIRE_121[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_14_Im = _WIRE_121[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_15_Re = _WIRE_123[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_15_Im = _WIRE_123[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage0_bw32_io_in_valid =
    Permute_Streaming_N32_r2_w16_bitRfalse_bw64_io_out_valid; // @[FFTSRDesigns.scala 102:36]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_clock = clock;
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_reset = reset;
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_inv = io_in_inv; // @[FFTSRDesigns.scala 101:34]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 92:34]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_0_Re = _WIRE_143[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_0_Im = _WIRE_143[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_1_Re = _WIRE_145[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_1_Im = _WIRE_145[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_2_Re = _WIRE_147[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_2_Im = _WIRE_147[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_3_Re = _WIRE_149[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_3_Im = _WIRE_149[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_4_Re = _WIRE_151[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_4_Im = _WIRE_151[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_5_Re = _WIRE_153[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_5_Im = _WIRE_153[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_6_Re = _WIRE_155[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_6_Im = _WIRE_155[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_7_Re = _WIRE_157[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_7_Im = _WIRE_157[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_8_Re = _WIRE_159[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_8_Im = _WIRE_159[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_9_Re = _WIRE_161[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_9_Im = _WIRE_161[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_10_Re = _WIRE_163[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_10_Im = _WIRE_163[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_11_Re = _WIRE_165[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_11_Im = _WIRE_165[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_12_Re = _WIRE_167[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_12_Im = _WIRE_167[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_13_Re = _WIRE_169[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_13_Im = _WIRE_169[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_14_Re = _WIRE_171[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_14_Im = _WIRE_171[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_15_Re = _WIRE_173[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_15_Im = _WIRE_173[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage1_bw32_io_in_valid =
    Permute_Streaming_N32_r2_w16_bitRfalse_bw64_1_io_out_valid; // @[FFTSRDesigns.scala 102:36]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_clock = clock;
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_reset = reset;
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_inv = io_in_inv; // @[FFTSRDesigns.scala 101:34]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 92:34]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_0_Re = _WIRE_193[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_0_Im = _WIRE_193[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_1_Re = _WIRE_195[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_1_Im = _WIRE_195[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_2_Re = _WIRE_197[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_2_Im = _WIRE_197[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_3_Re = _WIRE_199[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_3_Im = _WIRE_199[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_4_Re = _WIRE_201[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_4_Im = _WIRE_201[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_5_Re = _WIRE_203[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_5_Im = _WIRE_203[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_6_Re = _WIRE_205[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_6_Im = _WIRE_205[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_7_Re = _WIRE_207[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_7_Im = _WIRE_207[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_8_Re = _WIRE_209[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_8_Im = _WIRE_209[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_9_Re = _WIRE_211[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_9_Im = _WIRE_211[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_10_Re = _WIRE_213[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_10_Im = _WIRE_213[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_11_Re = _WIRE_215[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_11_Im = _WIRE_215[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_12_Re = _WIRE_217[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_12_Im = _WIRE_217[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_13_Re = _WIRE_219[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_13_Im = _WIRE_219[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_14_Re = _WIRE_221[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_14_Im = _WIRE_221[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_15_Re = _WIRE_223[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_15_Im = _WIRE_223[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage2_bw32_io_in_valid =
    Permute_Streaming_N32_r2_w16_bitRfalse_bw64_2_io_out_valid; // @[FFTSRDesigns.scala 102:36]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_clock = clock;
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_reset = reset;
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_inv = io_in_inv; // @[FFTSRDesigns.scala 101:34]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_en = io_in_ready; // @[FFTSRDesigns.scala 92:34]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_0_Re = _WIRE_243[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_0_Im = _WIRE_243[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_1_Re = _WIRE_245[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_1_Im = _WIRE_245[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_2_Re = _WIRE_247[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_2_Im = _WIRE_247[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_3_Re = _WIRE_249[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_3_Im = _WIRE_249[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_4_Re = _WIRE_251[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_4_Im = _WIRE_251[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_5_Re = _WIRE_253[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_5_Im = _WIRE_253[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_6_Re = _WIRE_255[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_6_Im = _WIRE_255[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_7_Re = _WIRE_257[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_7_Im = _WIRE_257[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_8_Re = _WIRE_259[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_8_Im = _WIRE_259[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_9_Re = _WIRE_261[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_9_Im = _WIRE_261[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_10_Re = _WIRE_263[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_10_Im = _WIRE_263[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_11_Re = _WIRE_265[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_11_Im = _WIRE_265[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_12_Re = _WIRE_267[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_12_Im = _WIRE_267[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_13_Re = _WIRE_269[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_13_Im = _WIRE_269[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_14_Re = _WIRE_271[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_14_Im = _WIRE_271[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_15_Re = _WIRE_273[63:32]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_15_Im = _WIRE_273[31:0]; // @[FFTSRDesigns.scala 103:75]
  assign TwidMult_sr_Streaming_N32_r2_w16_stage3_bw32_io_in_valid =
    Permute_Streaming_N32_r2_w16_bitRfalse_bw64_3_io_out_valid; // @[FFTSRDesigns.scala 102:36]
endmodule
